PK   wH]Y��l��/  ��    cirkitFile.json��丱�_�Q��}�Hb���������a���՝{j*�de�e�@�2�LK*��3S�L�����1�����)
2x	�r����W�fۯ~������7��m�c}�W}{�~}��mV����ݼ�%��v?��U�����2+�C��
�UM��.ZU�e�Zk�@^۷+��7o�}{�r	Ė�W%p����� ��pJ�� ��˶C�}���
��s�ر�DϮϬ
�Z(دP0_��J�+��Z���P�_�+A��!0�h�U#��Q�G�������~�"kCےV��J�B�U��L[��ژ�������yn�L�-��͏�Vm��]v�h�~sWo׻�c�nG�KC�#�}�w�r��6[D�p,�$8����F�v�-"R�R��H�o�"tj��Q���u�Z�߁�"��!3P�7�l:���ܘ�����H�oA�""�e�^�e6�F(��a���eF*��8�7�Flc\�s� �� ��nK�$ .��
�J�ey��Mt��?��o�-�ef�����r#=��,`|�;@�V��V�r�x���o�-w��;&d�q���r��,�`y���_���-"R�R��r�֋-"R�[/��H�kz�2��vǏ2�e6��!Gq?bu��F�;�G9�-c���ֈ-"R����H�o�""�E`��+�o�""�E`���x�-"R�c��H��"�""`��wz��d��|��)���-"R�}'[�^|��)���-"R�}�D��.��*����牛��`���,��E��	�z(a���`ug�����N�,Vw�;(a�b�՝��JGX�����cu�#,]�,`uW`u�#,�^�XݕX�A�K�WVwVwP:���U��.`u�#,]Z���,����z����:� �0N�׳�bL�X2x�v�? V?8H����x�D�P�5�1�ף3��T8�!p���#0_�`�8����/m���`�̗6����{�|�K����>X>��L��mp��#0_چ�8����/m�=���`ϰp�b�����|ǻ� ���/�`�/�כ�d���Egi�!�������|ɾ��G?X>󥭘`���,���&R�������|z�})��	����<Yp�d�����|i�,X��	�G`>}���?p����'f��NY��6��6�7p�e����q���/m���`�̗6����~�|�K���G?X>���`���,��Ҷ}�������|�{�!K�'�g��q��`_�μS]��ǁ�,�������~�|t���Kf�����G>S����z!�� �� �Ơ	��\��c.��8����/�:�sa�̗�������|�K�e���\X>��8`��c.,��RJ��<x��G`����?pЄ�#0_J��8h���/%���`�̗RW��_�|�KI���C�6@'7 �xp���#0_Jt�8����/�h�`�̗�ˁ��?�|�Ki��+�����|)�X���G`����?p���+|�"l�CJ�wm�5FUM3�B[7Uk3=�za��D���f�\X�4�����j?M4���i�؅�OS�.,~��ua��d�K͆kvL�#��M��\Z�iz�c0��g���ɥ��79�q��a���ĥ��79piy��M�[Z�i��斖gڟa���H����79�kiy��MάZZ~����T��H��rA[U�����5U���������*>�����CShWU�;��YW�Q��mWw=Y__x�����U|�ݳ�3�}�첊�[]ֺ�y�g��|��̴h���t�}:q�>_�Yř�>��e��c��t����+ט('SI3^��e��:��T�PQP�iQ멮.}LY�/���\xN�y7�U��9w�/J��Z{�J�T�Tՠ벶V�e?�Q���(>����z�i�����zPn�Xҗ��}S7�"���xGN��^we��*vYB���Xq%);�}?]�R�#����]���t�2���-�j��T��cٲ+��R˟U�B��]�w}������;��J�u߄�5z��9�ǧ�:�_�6�vs��޼���m�ND7�����,	J�FAEe;���FAàM�xD&	jMՆ�y�s�:~�<"���'A�Z�K��җ�I�Pv�Q:z4��
Q�d�l�(�'A��b�B��4̋!z���F�8r�A�K��Ֆ�D0�QR���f�L����L�$���rL&��FI�9Cގ�$A�`�%I�3 &�$=�B��@��8�b�P�
����$~���8J�gu@L��cI����	����ғ$D{g`~%iL�	j�̏�GI��!��JO��=1=�:b�t(Iz����0?na~%I�3� &X��R,j�����^0M��� &��ǟ%���,̏�%�S#lT����(I)��	%)e��1���y_z�a��~����nP6��`~%)%��1�����Q�RR̏;�GIJ��aS?0?�a~%)m2�1������Q��fhnv7�	����Q��FX̏{�GIJ6aL0?^��8JR�Xc������$-�@x��.u����JgX�qK*�U�N��¥�*�J"�zu�?.�W	VaիӼ9p�@�J��k��D�z�U�	Va�� ��f��h@��DXcED��Yx0�`%V�:���
ԫ+����i��T�^%XI�U�N�����*�J"�iM�L` q�ВmZ�,�[��K(쒉�H&�"��K����NgW_����d�/Z��Mk�et;�j��@2�t��� �d�0Z��M{dt+��Вmڋ!�[�hL��dhӞ��Dd"�$C�����V&*�%ڴ�GfbA&.�%ڴWIF�2q�-�Ц=W2�����32q����DhI�6큓ѭL\&BK2�i/��ne�2Z��M{et+��Вm�[)�[��L��dh�Q���e"�$C�����V&.;C�XF'B����,L���DhI�6�=�ѭL\&BK2�i��ne�2Z:G���Z�ŊB���+��eV&.�2+EhI�6�͗ѭL\&BK2�)ǀ�ne�2Z��M�dt+��Вm�� �[��L��dhS�
���e"�$C�rp���M#���-���(A&.s2q�-���&�����Dh��l���3P������"��DhS��
�$��Bt+�9�����e"�$C�r��V&.�%ڔ�HF�2q�-�ЦN2����DhI�6墒ѭL\&BK2�)���n��|�-�Ц�`2����DhI�6�8�ѭL\&BK2�)W��ne�2Z��M9�dt+��Вmʝ'�[�,Bi>d�2/�y��L��dhS.C���e"�$C�r2��V&.�%ڔ[RF�2q�-�Ц�"�-d�2Z��M�>et+��Вm�Y*�[��L���hN��a�C���m��ƨ�iBh�jmcf�a^(e&7�B)3�dJ���P�L��Rfre/�2��z���|���d�^(e&��R�/�z	c�s�.�1��P�����ܙ�K�`�x�Х^c�s'q.���S*���X��Y�K�`�x��ťb0Vl0V<w�R1+�;:p���зT�U+n{Sծ"���mUezR��.P�T������\��,)W�)K��Z�CShWU��ש�]W�Q��mWw=Y__�K���zɒrU/YR0z�j�YR��.Yږ�
mWƚn�j���i�R�A�V��(K��:ʒ2��0���)c�j�aH�ZGYR0ut��̒2���ՠ�̜#|�_|]v�q��M�\A�
�6���*�겤\��9R�{�)W=C����\_�^��ʕΩ�m��A�em�.ʬo:CJ�7�!�v��\�5��u�w���A��� _��Ma�`�����)��Rwe��*�:B���X�%);�}?].�ϐ%�*���P��S��ؒ��UMQ�JuQv�Pe��YR����}�ת꺨ݺ3��tP�P�M\���gȑr���(f�۬v���y��G�ˏzJ|���n[��-?�	$H��
!	��7!	ң������C�@���W����!	�c
B����$H�#�"� ��ƸH��ƹm��&��FI���{�w�y�$����	�	��Q��~����s�(Iz?�a��q��(Iz?I�a���qp�70?����sa&�70?�����t&�70?�����&�70?����3��p��-̏�$���+�	7��J��q��(Iz?��a��q��(I)W�	��-̏�$��T0&�w0?���r!��`~���8JRʽc���a~���8JRʑc��q��(I)'�	��̏�$�����0?���r��`~���8JR��c��n�7a~���8JRڋc��q��(Ii�+�	���GIJ{-aL0?^�������&'�r�R��RI��DX�j�'-�W	Vaի�~\�T�^%XI�U�&9��R�z�`%�w��u�	�	Va�� �NR#A4 �J"���"��IZ$�$XI�U�&9��R�z�`%V���CBK�U��DX�j�	-�W	VaMk�e��K��dh��f�
E]Ba�L�E2��D^"�$C�֚��V&��%ڴf^F�2�-�Ц��2����DhI�6�a�ѭL$&BK2�i/��ne�1Z��M{Jdt+��Вm�#�[��L��dh�����L��dh�^%���e"�$C��\��VhFLhJL&.32q����DhI�6큓ѭL\&BK2�i/��ne�2Z��M{et+��Вm�[)�[��L��dh�Q���e"�$C�����V&.�%ڴgWfa�L\&BK2�iﱌne�2Z��M{�et+��Вm�.�[�ՊB�e�2+�Y��L��dh��|���e"�$C�r��V&.�%ڔ+AF�2q�-�Ц�2����DhI�6宐ѭL\&BK2�)��n�L\&BK2�)���ne�2Z��M9Qdt+��Вm��"�[��L��dhS��
�$�J&�9�����e"�$C�r��V&.�%ڔ�HF�2q�-�ЦN2����DhI�6墒ѭL\&BK2�)���n�L\&BK2�)7��ne�2Z��M9�dt+��Вm��&�[��L��dhS�9���e"�$C�r���V(ˇP������e^&.�%ڔ�PF�2q�-�Ц��2����DhI�6喔ѭL\&BK2�)G��n��L��dhS�O���e"�$C�r���V&.��<ڃ㼫~�P��k[�1�j�A�ں�Zۘ�s�J��M�P�L6مRf�x/�2�y{���\���d�^(e&�B)3�J������@Ƌ�޹C_������ѪK�`,x� ӥb06<wL�R1+�;�s���X��)�K�`�x�,ȥb0V<w��R1+�;�pi�������u%0V<w��R1W���MU��TpZ+�U��I�κ@]SU����˒r����\��,)Wk�M�]T�C�_�Nv]�F�ʷ]��d}}]/YR��%K�U�dI����fI�j�dmh[�*�]k�ժi�?��K]mL[]��,)W�(K��:ʒr����\��,)�:��HfI��FfI��D��.��8��P��J���rM�ZOu�auYR�{�)�=f���V�%%��:��WE��r�s*x[�j�uY[��2�ΐ��MgH���3�\�5��u�w���A��� _��Ma�`�����)��Rwe��*�:B���X�%);�}?].�ϐ%�*���P��S��ؒ��UMQ�JuQv�Pe��YR����}�ת꺨ݺ3��tP�P�M\���gȑr���m�ϟ����lW�7�no~\o���������~��v���ͷ�~|���MuA�z��Z�����6���)۶�cOss�B//O����g%(� %S�3 �����-�肉C��s�c�k���3Mex��\�i������*��Sq<6�!qU��܎7p��>�5�%`z^.�u��<Y��������h2�gi2gk�4s�#�|���|9�����-\�Y�;���@�(�`Yĕe����I�0��2ۭ�-��^�������&��Y����\l�^D��/&���M��l`NӚqq�b�\a<�l��`<�>� ��6� �g' ���Y��i:	n��X<9�}���O缻eA�4�v;���&��X�vV;�.�i	.�yŷy��y�}�������}wn��ۈo���o?�����'~����Eq<����x��h�xR�0�	� �|~�.0�
��ϣb��t��/`V�Ev��)���SĐ��)>��/�bq���R,n��}֟,����c��D����	���X�� JG��A`�o�_����o?�~QK~0P�? *� `F��@}�W�{����'���`İ ����9̙�\��n\]	t�(1�j��K1T������@� �	?�rA�sD�J ������� x��p���z$�>��D�kw1T�%��J^A/������_��	��ϼj3�\<|��*���.d���q�}�e�_`�(�ZC�^4��B���	$�]vG��X�q}�Y=��]����a�?a�۬��͛_8�KYaV��-B�Ye���������=�[:���M$2;Ŗ_�v
��!�1�ֱ@3��5���[��k�O�kv	on�w>T1�bu���ݎ	UN��n��C�E�158�"L?7����2Nj�����\��W��e�}&���IyƯ�D�}�u���2�>S������p���|z�:��������lz����Q��m�:nn�o ��/C��s9�xjf?d����b����� _l؎��̂�jb5z~��ʹ'��M��fp�|z"Éz�Q�9�LOm�t�Y"	/2F� �͗��Rp9�2��D.ǙN4���ё3�#������q� �ޟ��Ś��G� ]l{�i`�qY�[��a�c�t��2"��͗�&m�|���2�I���,s����n�e�k����F����2"�5�eD�/�ˈ �˗9 Η/C�<���eD���ˈ�n2_F� ��2"�#̗9s� ���/#r �)_F� �S����|� {�t1�� ʗ�HpLd,_v�S	)o�:K�d'���O�x ����$�:�|��+֟��G`>��`�Y���|��X�?,��bw�?����|�[ �_����|zU��W����#0�^U`�U`�a�̧W�� ����|i=(��H���&L�W�:�G!�0�:9Mr�et(2%<��e��iY0Z���LHh��.N���bj �L��@�,��Y���&LK��:D�-`BB�e�h�c0!�	�~�����Єi�Z��LHhB}��3���b��Ӭ��WFG1ŀ		M�v��u�O�O��gT:l1�LHh��lg^	[43lOS�^��������b���&L���:DG1`BB�ch��0!�	�n7��Q��Єz�~*��	�I��7�j,:���LHh´��CtP&$4�>����!:�N��^�l�����׍���c��q,z���Єi/Z��(LHh´��Ct&$4a� ��!:��0��F�ŀ		M�v��u��b���&<N}�Y�=	
.�I_�00��j �8t&$4�>ʎ��!:�N���3��:M��W):���h�y0XO2�CbT:!<��̙ 0���r�
Ĩ�	S���1��Є)�Z��LHh4�Ct�&$4aJ���!:��0%��У�f���&L�v�:D5`BB�$Ah��0!�	S�#��Q��Є)9Z��LHhX
�C�^~�f~t���q�G�)`BB��^h��0!�	S22��q
��Є)�Z��8LHh����		M�ءu��S���&L���:D�)`B�F���][��ЇR�]�*G�QU�*���M��Ɯ9Esa�IŅ�'���$�]X~��ua�I�Յ�'�R��$8]X~��ta�IBѥ��6@���'�-�5��!rKp�pzl�R\C�����q-qz��R\K���T ��Gh-����)UKp-�p-qz(�R\K���T ���-p���T��H��rA[U�����5U��K=���� ���*�*����UAU>Ğf�n֕k��|��]O�ח�?�����*����s���f��`dmh[�*�]�ժi�?��K]mL[]�V���*��!�N�Uqj'�<�v.4SY�ϜM^0ĝ9�6��_�]c��tS(WP�BEA��D����h{Y�/����|_N��~V���չ�(�*j�+�S��RU����Z]�W�݌��݌���U�R�m��ީ����E}Y(�7�q�)Bh.�*䔿��uW�z�b���O]��+I١����bp�����*=���q6�����)�R颎�ˮ��mgV�Km�wE�����.��j*T7�}���_l�s�������r�n�۬����7���t�n�|{�VЧu�鼲��1m�N	2��K�Ij��OS��Y��6��m��4F�8�>c�1��qq��&t<ͤ&�0��I%L*aR	�J�T¦v�I%l*��o�ft������u�6��u��������s8�����c������@�wsT ��
Dc���}�K&�����VU�">�tr���ߓY�) qY�
�yH���E8���r��3L���='�8��zb�����L��'n.�k֥�?��O8M��Ra��)!�5��5�u��B�S�Yjg�x_�x�;���N��#�4��TC\f�M�in�)!�{X�)��Ƃ��:�;M`N�J.��n:����d���S�29�=�a�c{Z<*��O�eN鸖u|J���)׬���/��N�U���W|�����[槄�ލce@�n#�r{7L���a���ڭ�ꦿK1�-�a�?��W�Wwr������y�f����5;�枯��5�|�O��g�)���9��L9��� S��?��ψg��K��R�t��^��.U�K��R�j��Y4}=?��O����q��8�>�<k�L�o��o��7�o�H_}w�:0����Yݭv�I�-�.(��F�aЪ��N5�o��S�z�eV��}�We��������кm�wew�Z�Z]�fh[U�mU�h��,W�}.�_�lA�z��Z�\1UۦUV7e��}�����=�z_6�k��\2�.]Ɯ&xR?�&�wi���O�l7���nݧ��X�m�w��}��L(_S��w��5{K�^Qq>��WF��}��
m��/B=���ph���P��CЃmۢ�9 �[�}E�7���]}��e�j��l��(����t����������x�y�#�w������ۏ�l��f����k��\��Zn�RyZ�����_w��z�A+7�ھ����^SE�B����(֔��)��*��Q��*ꐢ���Q��tUc_YU�5n|ZE�����uT��>�Q�O�E��FG���57^��a�����=�˽D�7߿�O?�R����>����ߧ���ۛ����cc�x����M���w��|��(���P�=���C����a��������q��w�c���}}�8���q�o/=�����a��޽���{Le��N��*��L����t�ԁ�0�h��U�;�uک��F�}(�-�B�e�Y��x�g0��A�3����;�@�������r/2ǿ��^��<���`7}�
��G+�?���R�V�Xv�����{��C!�f����R���7w���'"?y�'��w}���j�}�����m�?�״�1�6��I������3&<�����}�o_�yx�U}�=\�;��������"��'���Q}F~�iK�}����J��T��>y����kiǆ/�͙�:�8ƾ���Fˌ���n�q��������>}	����Q��G��T4]Q����rb��&6>��P75�Bf+�1�ć�?~�Q9��z�����T��R�y����B�>�2}v"�!k�;����Z���Ke_�~��T{�Ӳ���f��ȵ�=�>&x��|Y0i��5�h�\��*F�T�&��%�ɚ��RCQ��:�ժB���4��)ǆ9����d(��J��;�V�Vδ��m1�Cٓn&P>�����7g��,���R�"k)X��Y�������nߵ�����~�(���8�����/���{��oS�TaK�|�4ut=��3�����������>%�pp����W��{x�$x0���}��9��<�R^q�W��}s���:��/w���E��^�̅j�D1W�ϕ�s%�)��mz���"�\(�Js%ܹUxV��O}s,궴�;��ww殓�lF�䮳�Nr?#lz�D�8эm�����뷷�|7���n�|w����}����w7�n��	M�l�+_�iۈ*�rU���e�?�����n}��}���l��"~Pm[��TӇB��7���v�e����*���=��-�P�U��b�2�zh�-������w���������p���=���mQ׍.�/����_�$�ߢN�{v������w݁�k�2�)��@+�D�7�F�`�!m��H����������)UW�Eշ*���UP�к؁,��j �H����?��0�m�
i���.*�J� C�Ӻ��QwO���?��]�>�;U�f���Wi������k��7��7���f,}x矞����7���w]�����zK�θ�a}ן����'�O���h8W�{�bgAաrc��.cӣ�y3u4��딵6ڕ��IݺR18�uCڄ����eմ�v*�Czf�Ů��Tۗ�0�f-V�!��h���+iPuS֪.t�����Q\��v��w7?l�ݫ�~������W�|����W��/���^��y�Jw�z�o��W�ͫ����MlT�Ļ�����m6��|_��ψ����z�ww?
ۓ���������V����O���У�14z]z��Z�-M�n��ț�c��$$>w���ͤ��ץ����v���_��{x׏��77!��z*��iɟ����.u����0��Ͷ��~�ۺ��Ď���j-��Xm���?����bg��f}�d�-{3��Έ��Eo��zW=<6*�={e��������~�M�{7ʎ6��M�����M��ױW�������/��0~^�^�A%�q{�6W��-�����䶷�F�M�؜�
��ʡ���i��CО�Jc��<�b�rGu;��J�˷�7���{�	��_���쿑��H�r����)<�^Zᎎj2�"����'����������Λ�0�ױ�S@�ǐ��r�r�A�'�4G����U�e>���O����ާ�z�J�|ʕ�>Փ��3N�|��B�����I���8�&=h�|����+��� U1��+�}B �0'�2�L >n���&0Ŝ����Ow�K���U���+�y��qGq�y�tNo;�>�O�oˍbB7`�����GY΋�nh�~e�z;�qG���۪ʜ7��Q��ێ���[���A�=���T�ڈ�/^hg�u9c@�����ɪ��]��_�	U.D�U	Q������V������A���6-xf�2�՟��皀H�b�!��T!�Q��sM /D��v�ZS�ۣԫK��$�M����aO�lf@���
��x`3�6��|_�x=��|�h5��k��Vz���-^إ<�8xw�q�Ǳj�m��Lw��v�y�Cݹ�_����M�X���qA���F�d����ovτ= �5 +g@$h@��Ω�̺y���BȚҙ�v�|��v�A/"����2���%�ǁzJ3vqr[Y̍�� Ȼ���B�IG)s�JFP�4�4 s���C�s�K��Pʵ����o�e*]m�-��P�K3�	6K�Z��"V�0�?_�e���R�����k��7�P�7h���-� (h0W;2/b�L1S�G�0���z���dz���ޥ)���]4��"Vd�r�ݨ���'c�g����rpw��R����a��=���~r��ZW���85�.�3�
�E�yx�Q�x��}�|�3�@��e�j�K_:�QAW�8����~��G�Ǜ1���H:Y��w�Ø1�J���ww�����u}����6�0���_}�o��c}�����w��i��o�ݽ�n�g����?�����M�7��_PK   �C]Y��<u� �� /   images/12ff1f2a-9049-4881-9421-35ee34297c1c.png @迉PNG

   IHDR  R     N]   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx���%Wv'v�<���j�n ���#f�`��� ��.cMh�
��B��U�"�bl���&��Xibl��9�3Ӱ�muuuy��L�߹�f�WU]��0x�^=�y���{������8�����g>|�R@�~�2N�h���{���|�G�{�vH��Q��D��
?EN�4'��>�7uc�߈�0�7C�D�i���[u:}�:��u�Ϭ��_�����@�I��F�Z�1� ������1z��I�]y~��}�����F��wǁ���F�|Y��<F��K�7��v~Ɵ��^�y�<�9?f��w�y>��]����J��̼Sҽd>����[�Rps2"k����Q=tA�Y]�����`�}G�D^�ɻ�
������?����0F)W�Ou��Q�{9�'� $���N��_���P�}��v�wH�<J拞4Cf���Ԛ$d}g�%�гs��*�v��O����	��~K&�a��N%���C?��!�9
<���?�  (6!?�����������s<��x��g8Lk�W"��gs<ƙ�n�Z#�]3�ܬWe���r�q�M��I��uX��t��,fܳ���4f�Hy�
�蓂��K7|�飰������1t�3 �pA�8D&Z�=}�C��n拋���la����:�K�ң�C����ǜ�.��y��J��v$���!�����i��tDt�@w�(���h�yr��3�(��P��;�4r�6�<�'��d&'�j��+d&��?/��� )8T�v�C�V��O=~/W�S�W��Қ�
,, ��k7�4��S�Č>��G�{���b�w�	+��8�w]���
K��u��}�6��"�n��kǼ#�\C��w�p�})�n�9��y8�s}����C���Q�9(	?��3A���}^``�R?k�بx�
��Z�OZ8>�$b7��w���(Q�lC��%�������
���aD�n��7��5`������OENlC�b�p�� 'qD��,�y��տP=�u��5�K�}�*��U&W���+>1c��������G��كс��s�Øb�ٌ��f�A�n�����P8�Q�ס~�Kao��B����?h�� �p�T�Re�ʣ#���X��5Cu��3�𿡲=��+��#�&"�3�n��ƏHX��m@���P����2�x�giZ��%�F�U�IT� P�w)U��D=�y���f����}�s�O��@ߊ�7����#�:������o���M��׏ r��&GR�ϙM�&�ǸNh]��q�Ó��a�q_[��Ԕ��X��
��Pg���P�}����\�<�U;�{����t���t��:�m�P�e�����ɯ]^ R8��!e�2'y-���̳~��zf�&��# �'v7k2ĶMd�m U  ���.?~]((�`���ɦ��l�\�S.�b�s�R(���8eRi��/��h6i����������63�H�x6B\���w~��Yq|��R@*�4dH�椐F/O�~��1�E���h��dz-����+��R �m0 ��~��#`@�\�d2�cN^��9c�����a)����)��r{\<pn|wd��B1���I����(3G�9�*�e�>n�=���M|��5L8��֗����������{��p ̂�4��_d��ө�^J�%@߫ݿz���>�y�|�v(��9����5ag�}Z���)�N�O&
A�ũ�|WHA$~c�O������{��P���L�E=~�o������n�[ Ds�My2���~��&x�帍�V����<�C����u0�� G�\��(��f)S����=p<��<<O��3��¹�I�����1�q5�4��2+LtP�
�5�E�c��dI�sG��{���/��n�+�=55N��iqa�f�u�R�,��|&���ڐjC�G�lF�v��ܧu�;������ݥ�W(}�R���b�"�w����3��"_�f�!�y-�?lv�{`̑D;��#���@���j./̐Ǩת��(�S��(F�)�/=)Vl�c�U�A�]W�������k_۾�#�Hy���=~-�cھ�Z��n���!�J5�0pL��CVy���1��5(���j_'�`r�M:�qj�I��ET(�����@�����`��� Q�H	ѾҮ� ������#1���ght�|��ƨY+PZ��Dp?�5�E��xY&$�s����G��^}�y:s��#�_Bt������&�ة�v���p�&�����ɢw\�LGY��0������I&�t4��?��4}]�}=a4��ȸj�D��Ð�4�-�$`!�8��G���e`��>MO����4MN����(�Y2FA�Z�:ml֨�hP�Z�f�ŏ�L�t*C�R��v�J,=�&&i���3���v�������]ʗ���P�����	������Y���D�^Y*�%}/!�F���F�DF�V@��� (����:U������O�k9$4+r-�����p"m���F�&7��B�\�ab��|����_��$B�܇�*�֍�ɜ/f��]�Y��d�#������:ֽ�L*�����@(8s���A��u��>ai��E�������y�0�>حCi�SNR!�&h��]���ׁ<W�v��=X�Z�ɨF��U߇�b�u` Tb��g��ӧNГ���c�.~���>�T���]�y����ʕ���� �FJUt�����H5���R7<h<����Q��Cj�1DG�����EFb�ċT�j򧄪�d:L���נ~�J#��=s��8y��fh|�B�F��^��>��zp�u�9�)��4��!<�n��I�z�������x�$M��Sit��:{�F�Jt��UZ^ۡ>�S.�v���Og�=>_�Ó&���h՞�i�{��Ởv8Y&2�U-�P3�HL@^_�[�9W3a��T��Cczfq���$C�cT;�"�0L�+<Z9L)i2�!�����$��R�o������0B ��ۺVKy����-b}�lC�ff`JY��۔��!sGZ0W�A�]���g�Uy���ïL�<�Y�J�Tl7�O��ZF�b<2<��^��k��g,�.�͉�(Ȑ~��n�lm
����D��B�'&�����\�Ӷk�����󥢚k܎f���5�B�/�b �S!����=��Z(+ܶ�*�s9�*�Xߛ&HN�_�C�4f ���n�;�EO���`�ٕ��2��,� ��@CQ���L��6*�=���H˵���z�>0��2K��p�hI�5�b�<��6K`����̠�T�����O�3O����25�����~Hwnޠ����):w���413E��<����Y���@Z�5�Z����]�z������W(����s�hva��:s�2�"�Y�3(7��(�Gd��m V��P�C�b�b>Ь��-�3���$G��'��8���P�'��R��(��!�c�Rh��ײ��U���j>�P����L �G�Ts'4�O��7jNb3�!x\u��@;�"��
7��ܟ=��(�u	�����M��m����Ϭq�6� Ç?G9�X��>�P3��~��+�Q��dA���.��}���?e��n�I�5�n����#s5���J�	�Ȉ�5���Bu.�Xc)������s[���Lu�A�I�vO�!Ś��]a��/�����=�.�ܙ=~x�HV
�ʒ-����!�Pl-Pc c�i�N�NBQ�~���������|[Y�f��:��V*kf�t.��8aGTuoM��ٳ'��3OR1�у�7���봼tW���<}��?��}������I�#���K����+�����ګ���F|�1�ZZ���Kt[�9�.��"���G��*�|�b�R|>8{D�
 BKU� ��c� ���N:�W� �:+v�G�$�,��o(P��Cu7m��X/56�3��9y:BA��2�z�(|M��f�d�(Β �ϩ��٫6ZꦀPr���Y�s˃r;:�ѧY���b��9�a�`���Xxh�-�p�s��Fu�5��/�'�_���z}�ieW�1�0	6u�h�Q|�9�*�Çc+�"m�?�g"3�t���J�zi4��J3���x���2����`U�
¢��&`_�#�'�O��x�Ľ�s��%q�� ����>�:&�$�\��؁A&�TL4��\2�Qk��@�o��d-��f�'�m�Y-��x�@g���ӧ����}�2}����c�{��iz���Y�?�j��R=W�#�7 �t$Z@�ˤh��st��)�q�6}��'��Ǧ��ܔ�v����L�\���� ���Z���&n0T�n��a]�I���F����J��	�:e��9���!G���Q"����7
����q�B�2	���T�(#hns�M#W�7f���-��Ƨ��(�Fɱ�(�B�����6��B�:A]���/9�k9�;�3<�G�-��~r"�)�(�I�����|'���&5B؄y������w���,�' �Y(�\�M��gh��'��n[<��}�5<�5�A����$�Y�C� pc ����x�������Ӌ�n�`#Y�!p�T0:���4܄�x�Qz�-*�Զ��*.P�rrP�2A��x����'��V���:�O2R7JB�H�k�����D=�8C�f���h�����?�Kʗ^}�.\x�N�8EiV���h�uT����D��\.Gs��R�&�F��ާkׯ����Dg�'���t��
նV)��S�T��!��u*i����Y�X��(9�>$ߦ�W���A-q�8�X~h'��10�WM�'Q�)��U�01M���h8�8yߘsK0}eG�#e
H��W���u��{r�t�(y8x�,�b������x�5�V�e]Tz�͆��t796�ک�f��t�{T.fh��e����<k�U}h�U3��ʓе<��L5�4��Y�"kW��^�-4��e�`�+�ts�hw�g�Q��Q�ӣ\y�����N��������jw:T,�Ŀ�Qw�8n�Ǘ�8���EB�U\�Q����(4L�HXK�:��)�Cf(�p5�(�-B9��dV�ZN*��uT�b�!��]�d\:13I�f�h�����;t���)����uz��<2F.�q�~F������>PRV�;���@��S4Q)�h�H�w�6�ݠ��g���3���AחV�4�P�8F���~V�wc6���M���6p�n�@b;�夋W�P7	)3�sEG��@F��E�C_ѓ���{1��g N=�qÊ���E3Cm��JB��]�;`
 �-J&GCXg��#{A�#B�~7ڇ�G	��?�T��{�ڬ�jLd�'��{���������L)�e�s�4�6��3��I�lψKE*M�ݦf�)6��HY�M&D��)����d���|�2F��� F�>�tE4�Bv������C�T�l����JDLl.���a}9�X�7c�S'Ԭ ԩ�N��@)b![���ʰmÊ\ͦ,�DGTG�[:�]���s�ն����t��Ic黻�BW>���M�~�W����k�.U��pˮ����%6Rؑ�g�B�]��1����'~jr�^�pA�񝟼G{�h��V�����&O��F��#/������Q]����HN�#�@&'W���6d��F�}�-�	���HT���Ô,���[{�E��̈́�i'#�^l��'1`���b'��V,��v���4Q&�_�Mk>��9���#q4RN,37����u�f���gH]?x@���a�������OY�*�ό6E=���n�����,���o��`@��f���f��BZ���$��%�0Y �ժ���+����┮7�h�ե��8��-�R�h��s>�9����E3����Q[���&�$~Cex�%��ƃ���ϲ ,�8�ɻ��vL���1�v��C�i�J_ud9!J��,ɣ/qj3�-�׬ѭ�W��jћ��N���/)ut���$����Dj�}P�P%l��G����
��.}�����`��{�,]��L��7����G��)�ׅ��*��SH���`�(@B��.\s���V�a$��M��kk�����5^��^2,7����1��O�  m��!I��ua}����+o��0-�'�JS�Ӎ���X��B����ciLsT��@�U�4S���h#�0;x�"V�S���+�Id�jc�6B�a�Dg��*�������*���7ߤ��r��]���������%v��A�cGR��Ǧi�R���w�٠��q*����u�֩�S4�/�'�hwm���+t��"ݿs��}\���6��NR��ȁ�#� N�,?���������Dq�%�
Qb*����Α
�:��|��%�t=LZߵ��p(��8@4�#�K�QNô��A�tX���"�P9{d�U<W�Kn<�"����(�瞜����2�%��G��[_{���[�Bٱ1-��]���ո��C����Ε�<���)���W_{�v[=Z~�N��Oѯ~�5j���m޻M��O�}g���/W� �9��d�īE�&-re���	S}�j0��l3��7})6i�'�ʬhon
,"��/4��!�oe#W2֕�
v�n�#c���c�!��)��J	ֱ��ҲM��$X^aM0$�ޣ���k:�Df�r��22H�ؘ�?���d�ܟ�}̈��C׶«h��k��R���P+5J�c� ��\��wҴts��ǧ�3O�ٳO���a�X�43�,3Ġ)�i���X���8A;[[tgy����8�!|S���ڡJ!G������W^���Iʦ����M#s}*p�Z�63ψ�����K#�f)�u�[g|�1�*��x>��0jT�@��!;Ir�X-�����Ӟ8uЙ�����f1P�)�!%o\f;$�RKih�*g�d������#�j��FJ�cK�4cI�c"�m*eB�(�ir</��������(=��y*OL� � 0%p6>��{��O
[��c�3�ܳ�����р����	:ŏ������A�ʌ��@ ]Oid���:�1&2�;��S��+߾]A*f�����S_��RU���d�b�;�s�\I�Z(q���յ�O�f�0~iS��J�c�����bs��٠Hl�� ٣f;x������Ֆ(���`���hFJ����D���Gdd�>}�8|ͼ%!Odh�ø6��!�J�j}�4�"�f��ijrJ����ML�����V�|V���5�S�ݤ����{T۫���U�՛���G�b�*���>��lK8T�������ۂ6���1j#-��U��|�A�A5�I\k�_�)g%�LC]�T��]�ɉ��\6�@��N�; �(�6ɀ�j!�J��44H��h$�TP$��&Gٷ�E�+�a.�����
�b�1o"��=
�?w�U�a���\����Ʀ�{����h�آb��3�yGxk?��������Tk����䉓����T�I��S���3*�A�֫9:(�M����1h�Лd0�Ѿs��@ڠ(�A��-L36+05��yb���7�I&�Kn�$(�l���}ZŁ�DsU�a�pTX���ahߔ�����S�����8Ň��rl0��6d�C=�8�����z�qR��ͤ�8���f��W����oT*����+N��g�R�R���LN���������T)U����s4�5^C�t��m�"�-K�'��1�`��5�2������ɺ�:��ޖ���Z�B�%t�s�ރ������{�n�w�e
�R6R=�tB7�'�$T�8$t^��"���
W�PZ*��O�VSd#p8RlEr��}-u=� �0	�	<�n�g�����svT^}�������w�ޥJ�BO=��0�D�s>�A� �O>�$�w�#�l=ZXX��Z������T��cfZ�D���=TE�b۲���8�@J1��$�0���=*�<P�P�$c�]��aΡ��ٽ�C�>pW1�04�,9Wd"	&��gq���Qmwb���E7� �g9)"l��f������$�l��^D<�0�(��ƻKVbr� �%�����&�YؤJ:&�L���~?�V�+��<������j���#.zw{G<�xO|�Q�N�#�����"bDQdU��(���1/)�+4���꿹ۢZ�&7��23��l"��<L���FH8���$�cy���I՞M`%��� ���az�R��%	���M /Kw���6��m�F�t���'��.2'$u�*l^4���UeV<W��Y�Rp�@Q/4�X�P��'��]ʥ��T,�X�ޢ;w��+��J��r�A�u��a��9?7O7nޥfw@���H�`U	�Ruq�@�R���h�Z�3�����{��"���=��=S	4�"��Vi��q����	M��� �H�V#�v�C���  i3%�j�I�@w���C�N��	.&i���s"��v&����Qr����C���:��� g\��8�Hk1�O@�0�X�Y [�:��<Ƽ.�e��6i��x=���M���s知ٙY^7�Z����
$��/.�����o���DeL��mooȵ��3���iff�R�4�߆�S��n�ɈTY��&{��[���=ֈRi%l-/ﰘ��(��h�9d)qg�;M)���G/ꋪ���v��^(�D�����K�,����)�zا+j $a������Z��甚��)ة+��>3()^̿�yB��YS�+��NΜ9�W�Q#ٿ�qq5 �0���4ݽ�&���b|Ϫ�CFمC��#T��ËW3&�vX5�"�^�D��I�<t�H������	�"]�bv*���R�)�w�.�٦��Zd#n�Pd����g��ІQ��{�Ist����\���v)��u��1�!p"L7)6+���z$U��_%!WQܝ	��mլ2�+Ӿ���3֑t���f�`�iV�oݿC���z�E+��ɤD���]ZY^���5����,�
EZ{�J��ܥV�#ׄy�ɪe�Dc��j7�26Ni�����KaGH@>����If��n�ʹ��vG����ѽ��u(�����f{���XM���o�I���&��"0��w:mV�;�_��b��EMDĐ���PԺF5 �����h�`,AS�^Ye3큁��53|���'(ß7��n����\�)�f���ooo3�c�dZ�o��Uv>���{@�����+*� HQ3�1��n$T	�@��3g#��d��_��m�3J�I�`HM�Hp*�~*_���8X/��c�ܧ4JRs�8��1��b�JWWʱ!K�zk=��+�tP;x�3�9�!�{j�D��K�������v �c���\C�z�s�0���:n�4c�:s"%�?MSn����8}�쌔���)����{��hgw���1�m�{��hocc��>O2���kW����dv�y�:��V���v/�+�Kg|���>0[��M�
]D��7"��
O��*r�J_���Z���o��w��<0:T�)�@2��(�r�!)d��)���ޞ8{��b&����L@�tj|J���
H�-93��2ܱT��C]G�� fb`m��+���g���j��n����R}o�fx�3���,`F���k>�J��&y��iV�KrO�*b҉��s���+�z�U�V�T=Pn���2�θ�*�Җغ"�mTW9�r��*3)��=.��n�xB��Y貪(Q%I��i��||)Hᨚ	�@������{��F�E�LX�P���G��T��j�;#U=>lâ.�"�!�����Y%��\��~�@��I:�b��i
t�*��k�#��#K�M�^�=#<x�Nd��V~���aS�&��+!��\V�液L����O.щ�h쟌өS'铏>��/�D��ϝ;'�E������U伽~��������?6O=h@���N-HY=��C��ۗ��<�z!��I�IC��ؤȱ�ٲ�~َ8D�9�Y�J���>ES3�T��)Ë+�NQ�;*` ����r�3��޾�uRg�wwoW�HHC��& _bFe��9%Ū��T�qS9�2���
0��l���6]�����=*�����,5w�b;�
&G¶��C���uF�2T��qf��y+�����1����F��!6drT�2�Sz:�u()�t��R$�I�uag_ň"�K�w�vK�"�AO�;��d��VaJ�� �ݶ�1͋��O_R�f�E�)��ض� ��kG���ᨺ�g��7	w�þ���ӌq�y���o�[�)�1t�����|#�mj�;doյm�U3=2,Z݀�&'	�C�l̅g�o�މcj�-���Ĝנ�c�+�tuW��:g0,���A��Y`���l�R��b$��}p�"}��Gb&��ڢ����Tx�M:q��>A�0�vs��ZbR���V�W�ި���2M�ZD����S��R��!�V�7�'����mI�&	V;�E�{I5��'~k�/�a��+0z-��W^�sϜ�V�/�w�R����Q1����<u����,Ts�7����G�$t)�E.b+y�K�x��=�Z��y�*�џ�?����~��V���� R*�؄99�$����_���P�=��-dhl|Lo�ҋ[��bqR�N6�U60m�Y��]�AlS�A<*l�}���vu����@��i(��I����鶤p5* Ir�+��P�3R�8��I�W,���B]N��ʨ02 �d[f� e�������P�G[�M�TE|8C���նX��ñ��ri�� 3Ô����]L\s�
mU�7��ጼPo�b�1[�g^�߫~$��ʶ��m���e��,�@,4����؟%~�Mچ��U���Ym�S�vd)�_n��[��m?y��k���_��ӧ��W_}��VV��K�*��x���]��o��k�ڏ��n�� �lWi�;�fmkD��1 ��n�<"�m��$�dne3)1uA�m���޾�L�C�)�F�A���3�1��*���1��HWx�����j=I�C�R<IӺ�z����&qxr�2��JmX{���9fu�"���t������~��l[�0�|u�$D�Y�p��h{�~}���d�%��D90��-��iQ��2�K!�cL�(6�C�� ���zq*`���^̡f�f�W�3������t�U�Sk�JޖJg)��+6�WBIR	�5�lJ1�N�.U@����뱶���Wq��	��m5s3��[Xjk��{ȹ2d'u��p<����J�	�&�������u�o~�\�[0�_��i*�D6kc�1[��6�0y���J� ��X ���T-���#��f�f�L��%���x��wD��@	RٷB
:+[�����р�*�;/O6y�d��		�˲�V|j4[t��%�S��SLf���Y��H1w7�֩V�3P�d�=�?����鉳��ŏ��˗@��q�}
���Y�רکQ���ﷹO:�lT.b@����B�G�<�q`cZ8#q��E��P���qz�1dD׋)�Fчc
�3�;�$��y�!,��y(�t�zL�U���G��g���I�Zc��P�;�fg v�N/�M��&�ٿxYg�y�T�zm;��Jg��#��h���ޘ�8|�P� 6�$��@�sWԼ.�{.�KZ\��,bQ�!g�Q�����Q�g���iku���רȪ��Ζ�f��R
�#���b���]-#%̓�v���xq������25�&`)]�Q���y�G���`e�G�����m�K���X����*jal�5�R�^N��w�#�b��k3ָ�������F��<��^g�X�r@�f�}B��
�mnl����G�hbr�v���+���̳����܌���ZN���Oh0wh$���z�Jսz�/Sy|���F����,-3��r��-�\ڤv}��,�{��qS������~��P=!����6m�5ibvB2%R3��:��U6�T1%9$�N��aY.�,�����$�`Lb������V�?%^�� *�i��E��ģz��j��.샑.�wty���0]������bu�Z�J�`�GQ��@Rh�e�խ��-q�Dz��H9��@/zɖ�qL.���١ '�&:�:�b�Jst��I����Z^Z���OI���	�� ��$�M,��R�Ǫ�`g�t�;w���1f`j����V* ���ؚ%�m��0���ð�o�S���e�b:���z H)���J*2�c�տ�=��ؤ.c�0� -���b��6�v���#E[$�%P�D]�9�X]�3te��x;he
�Z��m'��5��F8��qy�8F�Ͱ�a�\�f�P�'�&�X(�*���n�����h�M޸q�Ƙ�����N�0���v_4�Ty��Nӎ8�n\��ZV�N�<.N���]I����^D3'樘Y�r�%�p��T��w;4?3%�'����2��`��'��ϖ\�՟��A�֝����K���{e�U�42�A�*�ja�����"������pg�������m3L�)3�Ѝ��G�v���sg��ܸ8�P)&
Ӭ
�-)���^J6�sܮ��6_��o�J��1\u��;lx@���&mno�bS('VC1qTb�Ϫ��3��b�{iG����޵�bf#'tu�km�tUX@�	��`u��͎�0�MlmmU @��R�B!��vc�,ݡ��	���+�^�x�"��B?#�e�<� s�X`fV�I�=�1j�G;y���(�e/v�S��o �&�C�%��|O�֤�v�Eqcd� La+���#�,n����v��_���'�Tߋ��1��i�[ֶپ�9��x�����!&,)��Y�0`�����$�W�����O�UgM��G�¬��f3yj`:��Te�V�.������czzFҳ3�hux���� �ݝm���}�B7K�v$vyG����ʝ���[oп��K�c��Ӭݤ�֍k,(���h ���Q!�����l���ݭ5������$nSr�E�Au�>E�	���B��T�9LJċ�p_&��a�M�	��*�9RA�~�%��N����K����0�adE���&�X18\�Z�Q%=�I���#�>��\����C�`�"zass3�E�a	��;���&��g��mx�Y�z�T�;�/6R�mp��	�^�*�+����{���� �x���0���rz<�,���P��V���*��o~�~���I�fRT����j�r0�S[eD�A$ �J��Og�i�Ϣ��t98��%%m�v�M��߻!��	�=��Q;c��FqƩ�������5�p&�����v��rb�o+a�FU�˾o%'i��.8d>W}@�YJ1������ʒD�����p�Q�Z�08��k N$�{1y�h(o�ZF$�U;��H�� Wđn��h��&�m5hk�E��#������{�٧�9�<�E�v��_�*�䃽{��?�g�}��l2`*N_j����RR��7�}�T����k��V%z�P�ɯW2Ep��& v�T�L&��D�@�KŜtr��N��5
�X��J�'� ����$�ȶ���١�lY&���.K�V�t>oj��}�e��&�� �6�bWR�:��zKl�'�=�A���f��FS&|Z��`*A�mq�/����N�l!�R���/g ��!|�{ߡ�^U���8�wp��Oj��[V�_{�-̠�CZ��&�Q���6f�r��,t���:�����F�]6��^���'[L��C�6H������v͊���cҸ����k�Zl�V�f���N㜈p�0Sk
[�2G&�4�B\s׳jmƧ1�_m+�^w�0c[-����̭�+�����)���F30z�����nl�L�Ԣ�&ݻ{WT�'Ϝ��Ȑ��e�8lf��i�IG��5�F	A)� ���9��T)S����{�O�i�.~���E�����}��2Ԭ�P�Y�9�+1�Њ����D�w��?����h�a�y�y ��v�������M/����J0=�0�2I.1���&� ����sۄ�����*��6���9%5�"1�iZY�N�\��T�Vrו��g؋3P�U�+��N�H�u^�SY�G)��V�wifv^����	l*�'Kw;�Zw�~B�� ��04�_(f!��|1�m�zSl�˫۬�<�F�)��b*��%|�*�~"��]ʤ�EjP l@��re�\����4e"�2|e���\��H TiUVZ$Pd"C�,T���i5�Ц��-�:�+y�O;45������a�nH���������oml1�����D8���0�8�
MRsFه>E�kRj?���F�흒E����1�TÕ��֦
Y���	ӓT^d�V����q�5�B`��0��!T�3��a�Q��7[�$�������wz�J�q��<?�����$*���n������b'�&{�I�#BE>��xJ0��%�%b�5~��^L1��'T�ϙl���s�n_�&�Y��c�2���9���Kl�j~���1�ޕ)�1�r}>�`V����X�b�t@�y��~1yO�HM��w3R�:�i^�}����~�-j��Yx�a�gx00H��(Z���J4B�|�Rk���qEp/<���.���'/K�S�,9���^�ʖ('x�},$��6�N��4��u���S*LQ�٥�7o�������]Q��h�L����d�k\e�z��J�*�$Tm cK��P��%���&=Xۤ{�����[��4>1�̯H9/O��6��As��8B�#T����O��d�������Ӵ���ݮS���{�;��f(S��60㾏����ɸ�h�T#��=�R�l5����t��S��{<��R�0�E�-�5���P�x��,����.�.k ŬG�S��j����� ���?�x��4fP�Q�Y4�w�O�����9l�+�|M����9IX�)�G��Pe'QK��?Ps��z��C�}sv.�)Y�vŚӲ )��^��&�!A�� ns:v���hA[5���n��q���*h�|^E��q#����R� %Lp��^�S�^�?���pW�=؍a&���vvuzg?
}H��:$"��F�Ōjw�YUGTJU�
Mf9=���7��B8��k[ו�zz�ar�Q�i��װ�kA�}f:=%麒V���~B�vEZ9��o*1�)_"P!B1j����U:�8B���.]���Yeɓ˥��s�s�#�D��Z}l)Wt��Pu��o��Áؓ�m����y{����F���`��w�h�R���W�MΝ����8s��٠����-������ߢ)����&���E����2�m�+/�@��v�N>��@�K��O���_ߤ\1�� �ZE:�S���;�g����iIJ�8��	���~(Q%79��o��[4�@��W_��=ê��HM�x��w�G~���CDQt�� 5�gL �-�Z�o"�,�#٣U_ z�C���f���R����Yk;Ҡ�4H������@m� ���#ZA����QK�΁J���������3�2�G�We#5�8Bh\TXHR�����T�)U(���lQ6�5�v�JǠd�t��~C�=T��0��:5;-�\H	;0	O�K(���jI��E��u*���|͝�*�&sT)�h{�/�;������%��:��BR��-Yk`x�`��cH�X�M:9���5�so��,�W{x�*���	`!	��ՕZ|�9��[oб�A����c41Q�s�����e$6ɝ��t����3�N����� [ ��w?\�?�˿sG���B��枾S�K�����,Rjl��N"(�Cc@���1Y>$��ܻ�&��/6%�VHS�A]6M��ێ�`��=�x$ D������� L����㪥�q��/��2�(�%��)��6J���q'FQR۬{�w�&�X[t��Ww�I�iTq�HB���J���;٢]�T�G��b�z�0r�"�}U�:�@�ǏS6�Kٺ���� @���S�XA�-���b�P`,�=,:8��*��h��֝�t��
:^d��M��yA�v����Po�[,%��t�Z{-�lS��M�cf����TFdr�d��y�uz�Ü��}�Afj� ��ر� ���I�vt��V�Wiuc��(�̙�l�Q6HGE���.
s,���"kk�����q�D+�o,��x�.��-+(�K�I�R.Ǫw�@}xR��ft�ǘS�	"��W�
DS�N�җ�RoI�F�Z���St��Z����Ο�c��T�n�p��{��`�?et��?���?�ö]�.I�<�|c�xx;�GQn:(��}~�D��Ю�p`L5�Lj�:�:�'zT#c(��1�"�z�FKKK��֔	�Mx���دт�����.d��I���i�ao��lI;;Q��=Fa7������Q!N(�&,�2b3�d ��Zb���l6/���I�������l3�l�×��*��Ɯ��3 ꐮJ�Y!š�l�J��R�Y�;�ɑ�.�����.=w�����+7�q�{�����N%?9V1#q�8fG�D�C�ފP!	��LZX�ޥ�߽H?��2�bF���j�P:W��N�DQ���Qf�7��wD�So�h��>]Y�G7�_���o�F�QZ�ܥw��}������g�{��A�;&O+
C�@D��$'�l��L��wc3����d�������8U�3j���B�=ծ�w#�r���������4}�ю��s��c�-t�����{0�Q�4j��D�@�0:�\K9�(Qя�M�!��"��`U؛:�7&8�*g�����V<�!�Y_ϗL�z�j�$Bd�Y��d��{�DMLL����;6:�My�q`;�PjV"��4]��G[�'o�ܽK'�ŁQݫ�6B#�c>�#�]�{�m&�&����n��+e����{���;
�N�ă��ڊ����QO酮r��7��LР������tbq���ڮV%����H�$TU�1��l�j�����PVT&1$G��W�я/~H���E�u�6��S�-T�|�Umzjf�.~����ү�U+���[͆l*�`徼��Q���bнF}x�.��<���s4�lPmmev5�DwP���'�i߇���8&3G�
�m�@�`g���k���M�`Jb�ٙQ�}�@un��y�җ��E ��xt[�6)�:C�0Fg�>խ:F�ާ�%���b'~�̝���N�G���N�?ӡ����q�CQ���xv�R��8����*j��p�MNL}�7$�(��~����N�y+e]�����z�s�HVW�Y5��>~�`�
#u6��8�{�����;t���e�.���<M�.���H�� {!j6�vs4h�T�����Qy�X����	�b���*�ϐ�j���-���)�1VJS��G���E��=q��o��$�"b��)��}"	����P�3ʢ_�^�M������M7��N���dսQa�B�|I�abO�����Bp� L�x3�U�%I�_���l6#�����-=���������*\��O��Z�y����C��qk;b�Ҙ���ԎͶ/�S�̤2�:ǂE��MԗTM.�{.�"Aҧ=l ���a�:�G2Nw؈?�cJ
��b7��@p$�2��f��Efo,�P�5�ǎ��m���wx�O�3q\-���׋$yH�dPhv	|ۮ�;	�C�7L�'N�<��
+~F�l:#�d򙌨܈�3P� q�ົ�-}�Y��̜T{"I�Tv84UaN?F7n�bP]aշEN:O�Ss����%'Z���o`?�2����8t�<$�u�,�n��٧��X�F�\�Uܻ׷�g��?}�FKE�q�>�|� ;�8G�c r_R�{��f��=�z�ai��Na��~|������N�v���.��e���9�w���n։�ʛ�(�	��I�R_��#��P�Ta����]){����'Պ�����t�)֡���X���If�:UR& ϙ��C��)�
���5]��0�(Л����#ß,p8��`CY�=DI,')a�y&��MXx����֐-�H�]�Ϗ>d,��;�+�)����`�7q�M��}%�k��CN�Ė){��;��k\�ډߊe=���܊t&\��گG���g:"J>H�pg��'���0��^D�FS�Z*���IBͰZ�#�?@s����$I�Lt�o,pԻ\Y[���5��[��gOS&W�Z�AFlUZh$�7lf�#����������N�Ycql�������Ln*� ړLt0RѰ4v 5����%P�\*3�l�b��t��o��W�G���<Wn_�+����O,���ݼ��,z��?��p�����XUS.Mةkl:æt2�c'`�nJh�Ǘ���7hes�v�ڮ�D��MN���BU�܌re{�A�L�?3�Pr���읤w]tQ������ Z<���H�@�<v'`�e�x��b����k�I�7�
 ?�P5��9�=�j��/<Y�)o<��c�]D�ސ� P�Fh�X0�LGT&�v��>#ĕ}�uN}�.�\	���*���;j�>X��F����v�g��E�2mt>�����X���4�|���� xܔ�U��v��LFGG��s0w�c�.|��,�,���M�������ڈ2п	t����Ʊ�}�@��*�g�'t�P:�VeQb�W�ڇ�`�2d�aM�5&�u�Q��%f�@�&c7����1f�ځ#q�YMax��w��M]�cԿ8�]�i�2�˥E]T�#�A���F*�.�����g����W�3�A�KHI^�����nG�S�<�? ɍ"ǥ��*�l��|(����"���t�����3���H����2��#T�����mz���4Q�����qH�oަ��-��������T�	��.O�L��ʷRTLDž�|�Y�m����ll�?�o3��0I1sd�G��YHd����bA�H�,6^�t�sJ��5����n��宪*���@m�,,՗1�E���*�(���("�X����4l���@`��v�􃢬Pq0����G�5�_���B�1 #R�8��{��t���A�4::*��`�"(��.ͧM��F1cu�/�$�J��#���|�D��� +�I.@���Hk]�"�E�����ޡ�W��� �h��Ph1�VWv�"*(��툠��b�A���G���:�Y����[�F[�M�9`�ц,��z���ʴ�8/������?�M)ϝ;'{�5\]�^��sD���Cm���3���mq�K���jy�Ѧ�'O�W�xS��׮�N�.�, ç�$FS�����L���	�~��Y٠��5�C^6_�i��{x�x0���{As*��$Sm��v��tyrD�2��O�H1E��Uj�m���M���d��ҽ���g����5Kg�8M��(���\�v��1�$��6O��^.�pm��B`�vk-"�r��Z<��O�IV�G�af�j3��U������%�ԍem�Y Ul�|�( "�/�ʎ����@��rN +�\��"� N �)�[�S�����Vo�yB*�u����e"8��z� �j��uO�m��-&w�R��3<_r�{��[{2�|���g,d ����~��o����?�7�t�e�(����b�v>���l���MQ�ۂ���%�!cLk?��� R|���󕲘#��������v _�X��l�6�#)& e���/�j��o��|I��cV�?]�ִ)qԪ$ #[҄Ғ(�S����@;~����ߥ��9:��"�W�_v�����c
�#�z�!@j�+���@`KC,j����M�4]��O�E�t�
=XY�|�,�baC;u-�Tl�H�i��9�x�^z�e�z�O��Ғ68��Ӭ�#b5%�3���0#���P?0�IcQB�^[a�%\
�6"�+�2�Hg�ɖ��M�������enc@�s3����]���`}�Y�&/��<ZV�����/�|�Asmm�6X}�����N��)K�&�n������69l��
�$�ta�,�\v`lFV!��	������.e%o\o��d�n4Zr>�G�U��n�M����>�8����c��W|���B��~;j�뗦N����^�.��;������������h�!p�x��~�"�=��ײ�N, B�b����E	��zg<�8Ԗ٪���B����[Z����68�@�-+u�!)��D��p�"&��u�Ā�8ȿ���$���6�*� ]ܓ*̑�A鮪� �6U4����%u
B{�R�Tvi��*[��i�5Uq\K�ZŇ�V���������N�:%����$� t���
��/�S�a��O����ɗ
ԋ��[v��z�*z�T��^��P��MMNI�~g 5
�$a��Hš�m�$�a𝙙�,�Zw�ܧ��Y�;8��d $��AE@��mw�/�=�d�ɏ��I])�e�����h���lq��E���햊<�6�Ƅ��r��	���Vjc�"R��j0��X���RxO�\{(����T����X�t�������O$yߪ�
3@��c��p[]�ac^���'�:Cs��q��_Y�f�X(�̴�d���� ���.����#��ՅL'M�񙁦�sR��&a�~BeEEu���W�W�r��_�*�m^������i�@��x�0T��VgϞ��07O��bGL�osR��`�"�rՠ�`3%�Jb�%]��M�	�Ȕvt��e3W٣���+)�}�3e	�X[}@��-��?KSS��4�Ӱ�(
H�����sIe{=�0Kx����`JR�H%$T5�@�5�i��V-ahPX��H�A�ч8)�����xL�y`��mJn�}9t@�:��Yb�����繧<���Ě�S)�H69�y�g��\%+���
:��ϝ������]Q)Mft]�a�aU�?w��ᎫR@M��9髸I8N���Ȅ*&,a��� �r]K7.K������Ʌ)���gUsc]vK�j�h�hd�,��Ѭ3��Rel�� YP1W�]�ٖB+(�� \a)��,rˋ�ʕ���T�a S��SJ=�Que����xTbֿ��,Lw~�h_��[��x��������>]�vUj�BE����Mz饗D��Q�ff'�W��[�/O���[���E���	Ӓ������ωM�Z��T02���5�lS1;9B��D\{���W�ΰ�?"]@&��&|�5uq:�Y�����_�1/IȞ`���x�}����ߎ�o��<6�?��#���y?9�yM"�%P����kt��&$��-��8dHa��!_�̤e�p� o،a�@"X.P�F�?43%͞��*uRol�G�Ov��%�q��@2�J���%<�j��{4�;�}�E����X��ݘ ,ؖ�Q��*z$�h�/3c^@ij����Y,W$s��rm�f����$'�U;Z��Rx�\���T�3���V�?R�T����~��R	^�� ���?&��ƪ�3c#�����_�e:���xUD! �����з���e;�����0S�����O-f��B�}����A�ɟ�~�HRR==8��:)a�hsį���S�d��P�*LBO�ľl���fhm�c'N��H��cz�3�\���)y�Z(��ܣ+W/����7�7~�����i	�ﳸ�_��o�}���~���}���Ï��L	�ڸW ��"�����P^��e��4l�Z����}�Wޔ
Pio�Z t�G��|·���F[!�=B������/_�o}�[�=����S�����y�s����ɈI)i��a�U{coU뀴X57�g;���Z��BA��t��������ѕ+W$�燹�aᜮ�E`[�Se�5�<O?���/��onlҵ��ؤX�f��[�AdդH}�
���,�+���ʌ���[ܯ#b�"�����G���[�~v��G�DN�����$[��"h>�� ���;&��T��ORasaֆ��~����
�����k��ty���}A�Eţ����A&b�1u@������aQ��L��`}vf��+��]��{����?�&�L9qH��L����/�;��(��ct���H����/(�����H�;�ԑmWr���)N"L.4FRYns��gZ�7q�4�U1�Y�B�I��2 ����
Ls�N�;��kz�+��7ޠ��^}U��m�wV�ڭ	�:��/��	��q������?;���0�tZ��BŖp�@�Ă�*��D���f�$�Km�� }]�<�����}��~����[W�'�͂�E����=�����Ǿ.� ]_���SO��ĄԤDf@f�����k��#"H��(�>L(��m��]�}�Tu�P3-7ގۄ'��D��V��a渟���}���-�]p��������H���я�֭��ƃ��qy��1����ԘԼm4bӞ��pG(#� ΄���4f[j���2&�ȊJ0Qp�!-f�9�?�?��?�?��?�۷�R�P��fua��iw�퀆�ZiB�H�I��]��5�7�kJS�ʹ�����>ʃYgIN���쓢�#�	A��@9��K�RHY��pp�����^��L��V��/c����s��@�~��<V��t�+��ǎ�����m�߱�}�Amfr���Ϫ�?5KY�Mo�ݟӛ/?K����izL�h�A�[�Pe$K�<3�J�ӧy`����\�F.��O����8_/O||�����<��ק2Eɓ��b�iC��"��ŋ��Y؄�����@2�r��e���P�J傪H�7R��eԯ~�w��7������|��t��Y���/~�!���{���it������F��>q�%y�:�*�mWv3x�^��X���rqL�����z�q�\"�ގ޻hX5���Y�m�}Ww�ik�N�O��4�8���"v煩2��!���U�"4{�د6��H�+,\0$�y�N�L�W�&&'E��0����Э�w�~�Ё&�?�o�x2N����l�{I*�])ߨ��gʷ���*(]m��C(]l�vh��@�LFB6��C=��|�^��"=��Kv�" ��������-P��Z�\���Z��D^�#4�L�@��j���!�J��~��1q�qZ�|S���E��|��>:N���&�ٟ��+����8Hq�h���C�j ���lF<lZ���A��.�X���8���m�l2�$}q�e��Œ�F3��Tc��ڤ�#g���+�F0��ڡ�B�Ƀ	��nv���(%��W�3�ˈ��M{Y	B.�
�dZ�}*�����a{0A .�i{�5���ܙ_�csc��u���o�������گ�?��ƓrBXa6�H䫗.1�ޠ�����c�oؒ��k�(S���(���40�����%-Ti����udH6C(��f>��,���;T��]��G�X�����]��D^�CQ�s�G�2��0=E/���n��ݛ������3,�.����rp�U��W�ai���Je�GR�@�<ʶ�`�*	A��j�TH�(�}���Ԟ������:Uw֩���}� ��<.B^rYq�|9���������:��{ TY�A���O�a���� vg+Z�f����dzi�h����x�eѨ�x�R	�G9I]��0]�$u�$�<��2��h�ŶF���s�b�y��=ګUigwO�5e�}�B켻��Cu`��P(�ܕ�D{�j/&�TAp@�V*��w�uEs��{�ᚭ��=�������*�ᇗx~�$�o0h���0��I��ee徼�����H�#J|��A�r6�BF��r�����]��ˉ����t{�����jo���bt�;/lM�	�Q������6�o?���eYj-t����fe\�וd���h�
<8e Z�R\���Q�?��+y������"���9e�\YYa��G��{�Q���ʃ�R�^�@��t����]����(�Y=� ^PY�)�Óf�Wv��@m��U��WoQ��p��lf�٨j��'��X$ V�Q0�VC"揟���)j���Fpx�Ff��s3 ��U��Yu�PЭ��I����!��vڊX����w�&h���>
uS�M�j���� NE�r��Z�͍<vM��f|,/a~V΁�(���.!C!Bt�j��!��s8U�Wi�*��{g@{	`�2��V��|W���0{��a��X�Q�q�g���Y��(#S�Sղ���(f�&NUT�˨�#�$'�+�☼{o����;���|  }��?���>�k c	Re-�@d�H@��a����=�$;�,��^�,�M�j� ڠ��! :���r��Yr���*�)���	�F����Z���L�c�A� <a���h��]]޻�����9���
 �"v�@>���UY��|ߵ瞣Q��ĸ\�z���C������IB��[F�n�ȥ�]��{5�u��V�Wy/yb?���X7czfH����p$����KH=���۲���x�h4��~��(��;w�R�fSAh�7b����t\j����X���ԜT5:k��mн�?/������g�")h�[*v�`a"2�=���3�A���0�_iTI����28<LJ?}�2:z���?x�Q��Ѕx[Ν;+׮\���q�q�"��'�|��zCcc�r���ޭ�[VK�2�h������#n7F�@l����H�ࡁ_��B�Vsʷ����T6%j�p����,�g�M��nF���#ޥ�)��Z�X,�g����C�]M���K�U(g�=*�R��ky�=�0�Z��V�R��筆 �Y�i�A�{��c7��黏�X��X���V\�|�^�� Ϛ���(�爛�e�Z��W�+D��B��G�p5W��%��^�N�b�g<í��-�Q�'�	���b�䐕>��ⴒ�&��k���6��:5m���ٷ�������;�����,�wNE������ZAΜ9+�����7\�e�bMע��zYʈ�����u���k7/�WpA`�p���Om�n^`e����#�h1�Ư��];\�ޫ{��68"�/g`KP�$�bMJkBZ�Վ�K��Ư�052Ya]��N�2�)��5��lmt觷�N��-^_��`Y����27*�i<��RL�<.@�ݽj4��ˌ|alM��~�to���5��iff���X����e����g����Q�z������ӛc���c�t�t1"][[���SjKjRP'!m~N���/��a��*�k�3E����|L:�L��!��#�<5�+�6yҺ ���k�\�h4��2ܻRaI%�������uWt�[�SUgU�D����ۦ15���!���H�$�T�޸t&�N�b&�n������ݺ$����fvzF�}V�:;�}.,����	�*�okzf���f�cW��q�u��M}stT#�6��#��AZ�Qg���p[��Tj4��C�4�&|�#�f��}�N�V:<��LV���S��*#i`H����0��%��� ���p\3��|;��5�ڐ95�K�}a/�wa@���(S�:��:nq�bSm�_���e�����)����F��J9����"�����c M����V�=:�Ӧ 3g�qd�VK{'�E�vtu�˫W\����>P��s4�������F����ΉlF4+�>ɘH-�:�庴jZ���Yч@>N�
��	���L�\V�;;��i�h����f��O��\N�<)��Ξ�}��Ѐz�a��Q��];�_���w�}�S+u��K��}������d����K��6t��Yg�6��yb}m]=/خ*e�
ձ zͪ��YF���r\O�WS-�a_�p^7Ԁ��vɴ�Uk��HN��!e��w�!t#$������75v��3S��hN/��A&Eׇ7�F(��]+�X_�"��V��u�� �nC�&UYGT���1����<�������UM�0��� vt��H@-�����;�w���b�E��=\H�����0>x��[+T���Ss�3�u�"����P�;#;���s�&�X�{���}�7�|�sŏ`��4� �GceU���5V��0��s�jee64�p^����7l
kѺ�^�z��uu�hy '�W#�#ؐ��M,֨/��j+4��N0Yn�7j�ޡ�gX��{k[+�����8���������uCt�2�L��ٵ�*{���b�iyu]�k���*Xv�M&���RB��%�Z�kL��0N45~5�Y,�M#~�Qd���tW`�4�Y���)�#���ϑ#���	9x`�|��X7~A~��O�����#��������o~]�Vj������-nH����F����\YW�V��.�lV��tFʄ��v�S�cff��D�k20<�.#K����+zmEҙ��=��xU�����Y�&��6%l�dv�,LMH_O��<qR#߻YgZZ^�b)�Y�U:�F�W���4�0��ƀul��Q�@ĞӨ�c�,Cu�D���*ù��ұ[�Y#]XXd����&-}C e����G4�i�6g�=5�p�=z� @���Ȉ~�ܸ(��hN�lv�m��`�[�JM�������o�w�n8��G���Z͉H:�>F3��cni�`��@�	cx�#�3:ɨ��[��K�n�㌭4'�,�n4>?��2����Vs;l�pO�$�~cI��`F֥A�� wB$
b�)��D<�+h$���?�q��l`"$��h�5R��ܥְ�C�S��ҵ!����b�LI82b<|<�4��BR�a>��B�&ݣ�"�`.���L�N�>�)�Q�Nޖ�c�]��� a ���("�m��IJ����_�����r��)ٹ{PlR>���d�z�G��S5�.P[jǐ��5%��k4�=���9xZ�WE���ߓ����z�@��*P߂�P�PADVXe�h׮;���?���y����/H��H�׮����{y���7�j�ik��"m�%H�V*�lc��ƭ-�Hg�e��U�3�)O|�3%�r��a���H�.X�|�+K���W4�,����Ȥ�,<H���&��� ��kׯ�Ɔ��$F��#�J�`vMv���Y���N0����{��ZAmω��4��D�J��rĮ;n:��Db52���o����\�~�ׂ���#�e����n���ÇhL7���аєJ6�N�iDS]�97�N9� h<F2�k9J:դ���0��xݪS�������4z�5�p�[6���� �	�� "����9��o|�}�9�Гɩn��b�DC��kM��~��p�j0599�렕���α�C�E���/	����h�����a]��ՕD�b�i��U�&��uE�ߘ�O�Oӡ.��F@-�IМ�	]N���c�x�
��6L*5<0&-��%�k#93�2�:?3��mLc�tw�c|�}�Lx�0��uB?J�lwg+�����r@������&�=L�`�� ��LO0�����y!e���{Y/�ՋF㱴�v���eɴ��1'Q�A���6��d�t��)5Mok��~~�Fغyk�?~R��5��-��O�$#�z��ݧ�g���߾(}j�v��%�=����%F��mj��y�iT�����r��c�o���˩�G���KĖ��$>����r��rA����M���θ��=d�j
��߿�i�@�4ݑ�b������6�+�5�cm5T<��S����E����G=�!���F�р�sS�����k��9n�m]�h#�X�5��p�(wtt���o���F#�Ȱ@�r� i���������d�䞻ל�w�+D�I�1����1K!��!Z�{��#�Qp���@�g���j�I�?j����a�6��$"q��^��-6pm:+�I�SI��u$ؼ�M���2�MxEM��KՊ�%nj�r���q}���/��h����b�w@��}���l*&�.0����&�^N7KES�j�$v���)Y��Q/��� zD#
`*&z y sS��u�uh���lNΫ'���WF:��a;�:IW�Xgmh�Җ'�"Җ��Iٳw�F�9�0��XaFP��կ|�Hz�1M�w2%.i����<#o�����}rTS{�g�<H�Pk,�I��U)�۪4J���Y���+^<Aq¸��z�����|������%�hӍ6�O�%ɆUy���起����d�֘�-M���M��FތȽ�'A��J&�I<�G��S��Gz@��Y�����\�zE��oH��f*��sI���_X����4����ܼH� ��̧?�n6�_�=�������!R���B������_����Z]Y��W���?�	n�jgCS�"'�8��t���m�ai�ω;�c�5#Q���csww��ᴾV�Tz�cй�>���ή֌k!�f��k���ﯮ�^���v2?)�u]wIH��� ���MKm���(4��Y��6O���p���U��d{ÏF_Kk�+"gN�Q��egHN>|�j?��2�K�]������ k
�G8�f�'�M��M�B��"���AC�����w �Z����u��}����� ̐&8m	�3����� 1����!e�2�6�..�+ ��^�Fu)�j�Y�Fa���j �E78��p��Ô��ݪ2��z[�)J����U|-p�,�N�Mk�����qY_�������/>��᪼�����3�=u��4o�9#Ͽ�<S����=v�	�f�E��[E��ˣr��IIVoؗ4�L%M�t�!D��Ш4,�t�tH�X�o������7�=~��(���.hT<$�Fv�}��	�.2��	6Y��.��:?'�m9i�k��͂����Ro>�s���p^.^�$YNO��3���h����d<����kL�/���H�\U'S��{�嗩hp�� ���(˚������XQGtF�'�3@^��?��>�3{_���@B���^��ؐ�-L���"�vU*D�`�R+ ��@�谮a$`Y�zO�5I�ԊAA�� ʤj ��!Je�P+�qnPZ����n�a�`���z�`z\"���PVI%�2���C�Z'^�X�# �ǫ���9\I"�z�I��1�k�f��ގ���e� ��Y���9�mp_q�(�ƐD�bL��Zx?���iK�3�l�Ε��gBr���u���X,R���B��#J�q������ں�4��]|�/��-��0��i�PK����2ԽS=m��H������4���C��S���^����r��^������M�kr�=��0�Ac Z��c2�o/|�@/�,xxu�������dzfA�v핊F�2�'�(�����F-QA�-9���k��591.����/�K5���:��D�ܧ�
P���l@�L8�d�"y�_���o˳?xV�]�,������tw����������<���r���5d� /���Ј$��+�iظ��ki�Y���\�~�F��>�y���p�w��2<�S�������st^]ݝjH����O���M��Vaԅ��'�@�f�����!��R��⋑f�p�0BB�"}ik�!�Ej��>��YJ��d�њu��?×7@����q�q$�)=�7�Fi�im����H6r,���#���{16�?���ɐ���Ԝam��n��x3]��d2�\�%���cNS��YkV6�(��޵{k�s�Z���''O�-�]z^E���Ç�܈\����}����rج�����Z\#�5<���<�5�7n,�`����`�����]���c���)����e؟��&�_�\����i�qU�ji�n╅E��~��G�ĝ%���n��7/�p~�z�^��Z�HS���N#�uHZ�&t:�Rݘ�JiE�j� �'���l�7$mP�:�	FR-����5������N��],��� ���h�!�0�%		൧�����I]�y9w���W�Q&�eǎ~��떁�ݲ7����r�0�M7絳����iJ�۽Я�����UΟ;��<������CII��[._���	��J����O�d���'�t>�F��VlD�~ߴܮ#0�%�S�\�����
1�|@�p�h�V������J�56���\*o�[WF(��<��EHR�Q�R��0�!Xjm�V�F���aAY�ܠ��Fj��ܑ�N|�J6U��5��H����ZY@}��N� [��Fr���I�)�;�jP2��"�%K��ڄӶ�F���S����ل/d����z��z	5C��r�'�ʠ��ȇ��
3����H��H�W�����W�5c���C])��N��!6�c" X�����؂��QQO2�������]Y,�@^�ąF��UɥC�3D�
c\Xߐ��~�������7"p�8!�R����MV#�5Ft�ޕkӲ�0&5@;�� �,Q�Mx�\���kR^[�?��I����W��¹Wdf�e׮^5l�\���e��1j��������z�%�L%јHIk_J=�ٽ=��g}��3��k������}-��,�C�G��2���W�
�#d�MT,��)h@�Y J�v㶌O�ɫ�����5��IP{N%���#��XS>����t~�Ѓ���kB���(+dDos~g_w`z�_�֭���ޞ^Y�_h��-���	c��L��3oH�A�@��O�2ǳl��j�He�{�(j�2�H�����EYڌ�$�-����!"q7If\��1L�l�$K�@�X7s�84I�jQǽ�hf���]�S#��z9��O�OJLwm��G׈��,�Fv�RV�����$�VX���/�j��e��pF�!����ĥ'��#��ҞNHk*!��,�b�Pc���H����0�d �J;��`�g��o4��7��K�C��zc1���$d�fI�4m� b�T�$YF#`��(��=�����c!��/�s������GVtAC� s�����K�NwO��H�AM�����4��w��U��"����tP��\B*jLA0�1�"����<{V����r��A^{��g�k�F	��n\t|�)��q@�>ĉ��4-�R^vh����1��*��ݒo_��E��>I`��WUu�EAԎ�Ȣ�����0Yz�+WnЉ��+f�Vb��a�(f�/����-��g��`G>ʲ���Cn����f�ُnn!�p��Ⱍ5G�l�"�	�^��5��&A33[�i���%sh�����؍��M^R�����8���"3�k<�L���GؼA��/FI������D�bf�x^0�āV+|���n��sͦ��6F�@������k�#ꆴ�(�sPˍ7��'"vD�@w����+��*�/����^:�ley�C��`�ꢮ�N^V��I�!5 ��K��wR�8��IQfY=c�Fv�6M�4Z\�4��6M/��C4��u�@_�խF�|u���ش�lr�b�F[�Zoo��<�)$K�M��=v١�����܌z6̾k���y��M9�曄'A���,�ߺyS�~�;���s$����;	�n���� o"J�vI���D��}�� I)jDV�ؠFj�myM�29zC>���d����ƻ�9-'N��߼L��Y5������B��� �#{��L3�2���c������;eymY�o��ZA�t��j:���:�e5fEur�e�48��<�8*3
�M�����E��X�IΕɶI6��:�sp �T��c-�Z׌ ����v�o\��4�����@��Tx�%����r&h>�N� ;���?��3j�O�\��&4��R}�wg}Cǫ�RVc�QdzΑd��j�-zG�����T�׮�uc�B٬[�&l�r��[�MF��&0������a��O�>��.�{��q�lօ7*EQ���	�����b�������d���0�a�u��jS�=0�-�7;��'��:_���U���1SDÑ��G���]���K����,�C6t��k�u���$�4�qHM�Nn�/:�G�o�ɢc�is69t��xH{��v�J_W����-Yg���a�!մ�c�Ο<q@:;z��x��uB��9}R�������ô���N�����Y���.zOW�\�"�K3����]L](�h*XG%ft<�Y �ЇH�*	voI�� $@ۿ�C>����$����w����.���\�E���׸�����"�F���F
����@V)Ɍ�\\�J9 &7+��~��I8j���ʯW��C'o��)��Z��Q��V�Kf�TC׷J--L�`���S>�'_R���=6*��F��,V]���|�-�n��W�c�K��C̯b�
�/�^Oo?���쇎���2>>I� ��H���M��$�ek4,����~; 
�U>KD��x6ؑ/J�f�j�s�����Xi,��g��HH]�eCn��q*�|�>bnDN�'`/�X����K��#w�L��,0��SS�o��*�Qщ�Vy��m2���`)_[�>T�t�v3{ٽ{7��dL�����e�z�7H\ӧ����#���?w���XC`J�ͣ$�d��8��Om�6�s�5�_��&�0����I�ܽS���hp�W2�;ݠN4�FTHi5h�l�R��6M�G�yy��+U���yj닄d��:��mhH�8��x�u7�R��#��4JN�nf�%Nr1�w�i���Av��ey��Yr�h�<uR��t���9�
����.���V*��҄�3�RL{^�\��J='��e�X�d��L���5:�}������=��sϲd1�)|v�NF�XX�r=w`����K��-��05O�Y��:OM�5M�	�{!�����(X�G5�*9=v<����l6/�� X� ��{[��F���N/���y������Gd��03�� C�g�u�SWjqi�0ȘfC򱝓M&R�6&'r��d�S�,Y�,RO�z��B���=L� �r"�N���md]�kd5�§ڈU�}�k�?��r�.6^j7%A菩*�H4���p�h���e}ͤ�t�"@4�����)�:�&�oi!C��� ��a}m�{�k �������|!Qr��>:�z�٭o@��~�ٳ����뿖_xIZ�:X3u���/���F���bb�^W4!���^�����#�-��#p�aM�C�_��q$�?6NV��z���~���G���,���͐�*���B���Q�%r�To@�σ-p���8F�F� Y����6$�����6D>Ȁ���#j8v�f���u	u�];w�1O�QIa�ʋ+��_��E�t�C��e�4e�'2�#�T�l("�ixy�@�.iƫK�����Kr��9N-�+#Rx�'Ȟ�N&�f�fYx�8G�'�7b�H�$�Ɖ�`{9�M�:�	]'B?R�|3���0�t$ˇ�����P/F��d'����3��EEԕS����IVW�������J��Rj�l�$X�����@����B�b\���ܼ��s|&��L�aW$܈m�枑�n��<W4_�%n�)d
C
Ib`�9��6��A��ts\�	(�z��o=�����B�������Μ9õ��e/h���P~�����`�v�3��λ����d�I�"Bݓ0��8�������%]��a���D\���.�ʤ^��M�����<����H�)��Q�A���qHM�Zr�b]�#��$�'�B��EN�3`9�	W�Fԏ��8���|��'T�<z�����Y1�ūZz:�0��\�D��L"�f�lpĮu��λSj��ڹЧ�'Ո)9�	����jld�!vل�8�?7����nV�`���\Zzz:UNOM� E S?�}���&�\."blc+#��[���c�x��\|�$�+��ak����nrG6	4�S��50�5���,I�j����h�$56��|������0�q��]r��My������<.��nN������anӁ�Ľ�J�#h6�I���#����@������Úƞ7��L�Q_E�JS�<��2�黈�0��0�묃�D0�x��n��~Gn\�OC�Uek>�T�
�E�pԘ��G䐍�� �9�s:��7����>e��d�5�.����:�0Gt�'ԩ?������q��,�Ȟ�/]�	�	�����291%7n��@�7�Eὢ� ���@�E�H=�?�_��p�ߕ�[�Y	~�AMZͲ�F�4�ӛp��-��9"���C�IL�0�S��E;u�1�����L.<�0�d{#�RL�<FI�&�bS�,k��K2���z^��tY��͆I��$�p\�qU�8��Q�'d�r��M�����C�L��!J��a""hC�R!f������� :�tŀ��aT���H��I�(fqaV���2B�<��@������H��{j��Vޮ����&4Š;VNp`��J���G�Is(@J�9i��Cȥ:���7f~�-��2 %l���4�|`���>��l���P��Th�8��������0�Tk+���-}�ވԯ	���4�`�VV�X�3XP��Fsvv�h�];w���0k�8���0d�Fi���F]#��E5$� A)7���eOl�:�B�@�{���a�A��Qc��O9�*Lԯ(���ΊI6�R�1�WEF��pp"�C��я~D���	���a,/_�"W�]�ٙ9YZ]&#�|�TQ�D�
*Lk�+L�A�uvf��!8Ӻ�/G����#z����xl"����_��F/0(�^�`.���ٍ�츸O+f��5ԐFg�h�dM��u�����"�l2�� *�Yz��ӶeÜ�t�����0)-�@>��#r��!��	F�lKZd9���4����7F���ڊ�v�<��Èr<W�)iV��s�̙L�z�6�b�&\8�,�N�)aL�\� -c2���2p���r.��3�C����&��3gޔ�{��bQWDW<����a�I7f������#�	�77S*���50�^[:�[k�nl���՝$0l�$%v,A(`�ܦb�3�324���t*��� �KO�;�����ki3<?�ɯ�MnQP��� ���.��E�J3�cM�a���l�7�ϔ�Aa"hu���z5Umt�)"V�:2N_�۰��m�h��Z[�XT�k`���@"��M$Y�X$2+��H�}{L:(���Ӑ"Ϳz�ܼy�k~zf���7Go1����V����!M�ф¹�!"��� ��Y0��<P�08��c��ƾټ���ps-����k�č���LBn"��ǲz�ѫ7��3��Q�Ji���BP5�JP�oL��[Y��6QlJ��H*�7.���}����K�v��9 sS��ݑ������#Xb�&'��T����q -+;@2<7��p�E��|/����q5����NP��(r�?aSN�������n5��Ad��Fk�q�i��� {[{+ܭ[�͍�	�+ĦH��*J9'�Ԇ�2cZg�
��j$^�il#����(�9D$�x���#S��@%��~hL]p�4�湱��ڒ�Ԕ��lQH�i���)��{�N�)�gx�Am�����آ}8�j` ���s������Ⱂ�2���!47ҙ�dH�2�͸� [稿�4�0W L�Ʊ)%45���G��pH���5��F��a����>%(U��t_�/�[�q���ZI���ME}�	]{`�:�F��_��%����?��=�3b���>9vǝ���A�a������F��+�"0lP+D�`���Ն��Ck������o6m�:�oq��jI��p}@���(�ި�3/�\�$+u������ʔ�h���B��e�⇎]&rS�I�ey �OwbgYt��-��o@&�Geiyբc�Ys�_����(#@1�I��P{��Q��Y\3���F�U��
0"�N��	� �kl�'�Ի�3ԨZXX���EY��2��j�CDEWlXD,x�~���Q
��=sFN�<�I�V'��@#rj��@`�� i<iHQ�1�������E
��Y�R�1�j�5����ħ%��H�>h�rL��΋��D
��$�Æ��"�$��@\��m�����5��H��Ѓȁ�#�07md�{{��ç���~�(�n��?1�(C�I�������5 d�������{�� B��]/�5a}iGw�ut}�>���?���5x�ԍ
llѮȦ��3�?E��XG0�dNB�ڸ+j����X��#b^�4��ћ78���/}I>���c�[��&�{�k��q�?)�O��|�u����D�B:\�A7��=5��a �׺5��d��ڢ��3��wd��H��~�]x�zD~N295�=���#e,�M@J�Ƴ����,���dec�q�j�����ޚ.���BGZ�NY�����i�}l�������=�p�`��C��p|��қ�Lu+5nZ	�J�H�0�	�Hu��?�XeQ_\�,� K�!;䘢 ^����n>J��6K��?(?�AJ�ܸvChI���AB��Fˎ�ӞZ��	��Bg��� �N�C���H�a���XЈ@���N&	Kg3\�ccc����K''�f0�H �������N�Z+Ѐ�5�D]��۲{��7�[3���ٷ��St$9Ұ1Q�>��u��ۻW�tdh� ��D��Bi��SK4a8���QC$FmQ7f�B4������}|��t�3N��Ϯ3E�������@��!��H�"�)�F}��@y}��^!�Ei��QǱ���1�Ο�����G��~���Qa\��r58�5b/A]�$;U��˳�#�G����SI���]���\,�D��)�X���f�en��q��$�=j���F�uc0|�����\-x�(���zՐ��g{1���Nx��F=��
'v0* }`��|q|�i��T3�5ɞ��[78���=Z�8�T��72|�O%�BA������i E=������p��O�K�A,
�yD�+����4�PK�S�H TD���Z��r�Ʀ���R*���+t4���w줜E���Eb�>��C�w߈n�P�i�g�)c[c4��:������gFz?���?��hd1��1�ע�F�.���_���57a����"j�r��\�q�69"e@���R.�l�:���!��p�͛�2<�+��z�W���㌫�G����~�#v��X��Č���9���:�Wc�2	��Aw�h��h�x�%_��a|P��l�LP�lY�`Q�(�x�pߍ�)����l}��Ȍ_�4��2ཕҌh���i�$���0��as���^��Ѧ�e]��"�#�h�}�SO�'>���/� ?�ɳt ��� ��ڇ�a_y�d<|�y@M �(��zoҲ��������ܩ�ds��\�Is��%�D x<�;�&�]���<b�2�'���̻�?5��)@���a�dj�0��$jU���\��ƎfQU�����y�ʺ�JԕI1=�B�k�b���Y	�?�&NX�?v�8hI��VP��ZLCH̞�=������D*+S374
�)]j�0�YTǰV�Ծ�וj�lK�F�����mH2�o� 7��M$3�x�00���|�e�v,�>N>?> �C;��2�ѩ�~]�|Cߧ��zB�&7�.�3�rkl��&9�m��9ۯ�li�DD����RW�YgD ah�k�g���>0�_D���cN>��3�)�5���? ���O2Z@���~�!�Hvå�Dą���2�HK�:A]�ʤդ�7���w��dHz_ϟ;G� �I��𙧞�P�+?U�����bh�Df ]��0)^�p�$����w�E��hP���� X�o�ݦÚR�x���&l$��L���|�[�U�"gJ�N�iM�aP��env�� D�0@�����`��ڵ+�q���x�]c)+����|���eg���E֨D~��uٵk''�m"` ��!�3"x���]JBI��6�+�:����ORirfl��#;���nw�����i&�e�c-���q���-}�+7e�F:�b�M�˫KRY]���r�l�����A5<�����/:S�VT.Ʉ���%���� 2���e"�t�2�Ė�o5��PC�}���z�i�I���]�fp���d|jV�g���u:|��+�֥)��M��kuHW�n�����4���4�P<���v]T--�d�*�&����=�� ���\Ji�vcLF5ڹ>
��`YZ\�;�t�T����YrȲ#��nD�����pm��������?�M�-�v��^_�FTcjؖx~� szcN,�{�D�u�m����?�_>���QkS=��+n8\bM�U���禘���,!��F�E�9�$���s�tW�SMt���q��wحF9������K�5:B���G��������o
�!�G�#��c�b�����?�����@��x�t�O�H��FMOM^��8j���,AyF)4ŰA1y�W�ɤ\k��;��u���s4J8Í&�L��njj��x����'?A�P��W^}�%��=��p}��������KM�T�I|���5�)��+߰���@�l�d�/r��t���9�J��',(?���Ȇ��X�C��9*���h'�F$�Q�-���֗%Y]��nMw����M7u�E>M�5A�Z�CV�6d~iY�V(��]��fD�Xw"^$`��C�d�hl�r�cѼ�͚m6�0JG��&�:Ш]_/�9�Q�ɢ.B�ɬh*��K?�s��	�	Ҧ��U�J///�j������|A�5M���'�)ܢ� cZ-���^�jU~���2=��F�S�tc�w��0����zM�Ҧ���ܸ̂v]#�e�x]�؉'E�L;�j�	u�	�Ulp�����qa�G]$��k�8f�'uc�]�51G��p�Q���]j���;rg��ӈjd7�!O��d�_^�h�;�Sl��@����8�j���jʥ*eY ��N�}v��Ǩ��2�H�����H �� ��~{�8��]�r�$D�$-t����&7��~���0B�/�����R}�pO��w�F�`y.�Q�"�/��u`N��ک/35���_P;��թ�#�x���#\��giO�K���r��5��Y/���$��4�`���Q%C��㷙yX7&^�˧��2BkJli*q
+iܻ$a��� �6D�|$��_���x��hG��E�zxx�
�ulj6�6��������m7*�Қl�ޑr�����-a�B%Oj���-��mS��֭7,�^<Hg��d�j|��4*2�.��Ad��D�i=th���X���[nJ�5'�U�!���Β~�믿��@YӔxnqE�j$y����88��-�)��ׯ\�ǅ���\-Ʋ�>�P#�XK>����3��e]�3�_Nj���2��9K 6�QA8RS���١)�.9~�]ҥ~y� ������oR/
��~�<�� ̇ԯ����p����O�a[cG��E�)
0\ �
�F�xQڀ��<L������	
��<����pt�T۴�\43�:~��&s��K�p��?��?^7"T818<�:�Y����_#0�0�(�T)3��+a�T�j�`P�:cSw��8��`l4 S9�F�ᲃ/���Ѱ�ܹ��K@�����)�1����f5�G?�����K25=�fd]�wvuАn���d��D �� ��>����8wt��|�r��qF�?y�9s�,3d/ĥ6	�"�.6�uנ�3:�h Kku�Kod;��$k����&�K��xj�� C��g#�AY��/TVx�[R�c��������#Ɉ�Eﮃe9��a��x�hw_����-G�{eg[VJk�29vC7�"'����XS�6]�-|�z��t.!)��*`2*	���{h�$��CΣ�z�����Ō�/L{��=�� �ѧ���?|F~��+��������)i�����F!�ԗ��Fݐ*�Y]��N�:z�n����:�"���t��ں����PkjH���KU?{mi]^���������闁�]j|74
��<������˯ʩS')�|��%9t� �R3�za2`����=��F�]�N������Gsg���c��M'N>�� �I��#�ф��'�<��,Ҷ<	."��&
�܏={F��!�j	6��`�qS�Z�:�9�bd� �=��5�XG0�٬#C��)A�T���?�4c�:8�Cmf���}z⍞�>F�>��4�tE6������N�sD������Op�
�M�g�yF#�Q~���S�D��Y���=j(;i9���N��7�俟|�I�K�86?j�����Yr����l\��f��^��A�{ �9�<�vꆥ����K1;���ec�egp�\G^����b�!��<��}{8��kC4���rT�K�#6V�ͮ�F1��*z�2dڷgP��3,횢�޺*��/Iii��@�6�x��H�]���-���i$W���i*Ʋ��u�j���$)5�u��&\��(���L8��	�
7U�3¹lRN�<-�<���y���E'�9�[^��ߺ����F�C
W]7��⪤W��;�G�A��
k�\�IC�I2�E˺:�����diT����r�I�a�e�f��i�tCܖ5� �k
�'�Х�y�aQ�E=ncc��J�6�g�(����]j�g����Z^x�E�fOk$s��(PF��@OXLݞ!��p���2���*F�����?�8E:L. Q4����n7!��Y��@��^{�uF:���詧�:��>{�7H���7e<����`�#
2rǉ	cr���o^�����k�&����-ʛuNA����ޡ�Ƞ�tF	i�E�5v�1��t���sL�a��)?��'�G�;３%�����w���ڡ�,J,��ɏ�L�T ZP_Gě����A6��}��{�����@>޽{�P��,��d�G��)���UQ3�FlT�$3�db �4p]vÑ��7�Y�X�PҀCY'Dl������,a@����{bo�8D�]��#���
�_imMOs���E�ê�L����-�v߁C� :96H�`��p���6�ɱ��(W%�k
Tx��UJX-$��M�E�"�75#b�l�>024�`�KEt�y���qX��?!w��K�I]غp���P�z@#������;9J���������t՚ }�@��YӸFZ%d�5Wؽ�$s,w��i}����F�ռ�ZIӤ4���nw��_���R��FM�em-#w�}J�=�K�����yYQ#��-�7~ɟ�rA�]�h!o����n��<#.�f�8Ȇm�MRcl�*�.��9{E�6�2I��h�4���^&#���*���U�ԓ�b�ڽF�d#���,�?�A�c4G��Sǉ��Q�~�ۿ_B'J�����8�롛��t��$a�8JH����Fm&�Ǡ���Z?OO"����5���Q��Q��5�pPs�>fއw�/|�O�����o}��i���u֢;�ت�>U���Vb_��X�B�Ҽ:���O~�����'���>$��V�,4�f�C㼌��J$}M�X�y�IZ�F�0�F�j�^<�Q[������T=� �O���Np �7��x����k�k��
�$|�q�&�>���8�x`��4��iv;0�R�m��*7dX=���C���C
���0y�������`� ����X'IE&����[����.��҇��i�����!�(IZh<���9R���i�ylj��I�V�p��� C^�/|�s,Q��4��CX97"j�;�Θ9������W��=e����Lf�1��V�sIӨ�袀r���ҪF��┬.����#���h�ҩ�������{bkጾ������f�kr�ژ>��F��ڥw;7H1&fH�R֣ae?J���C�84���nm:Jk琌��� �%�q�!-� =L��%	�t�y��H��A{4��È���B�1��Ʈ}찣���z�!���׮IA������v������� ��5�{]ֈ��F�͌��W�����X2I��U$h�ppC:� am��j��y֡��O����6��'?�I��;�c{B������ߖ�/�Ys��1Y[_� �+J	���X6B���|�_���G���k_����ٟ��됝�����p��Pb�Zm����ҔR�tZ`��6ᤁQ>����$���Jb��4v����0�D�&J� �b���c�����c�ILJ�գ��3Dp�G��)67렱���xgD*��8����ْ��ּ�db��t����;�B�B�YP�Q��M�[��� o#=��S��%�Gǥ��C�hZ�g%բ�l����71��msČ	&$j(W�i\Z����v¡_�J�4�����,�	�9Bs0�(�~He��岃����"�a-�wQ]���`��4ZS�d�ٕ�>��F�����~X7�L�xˠF�s5���5�M�O�7����,����V
��a���3H�CT����9&��@k�`Ǿ��)+��2��'�9m����^6�I'��`@M׼Ψ��L2�VLx��q�����I��=��`�lڌ��'�І¯|��2zk����.^b����a��
5K�=
`��i�>gw�}D$]㋑�v :�1!�����}��,�<��g���{���c2���5k��ΝkB��(���D���u�>���RZ�3^����K/����1����YNV9B'���OQ�o��l\6�jB��zޡ���:�	�8���A�^��?�֔A�lSN�i�/���Ł�� �l�9v-�;v6���l����iH��bK��uwv�����R*��]w�+�������5m��)����j�.eG�2����O�]�F�*�ըf���eZ��(n��2/� ��P��7=5���E�p{����nRB:��e#v���)�D�5>5�)uI�w.�x�5LZ���p�]]x]4yАW+�V�h�S1���7<"'��)O�q<�h�`�iDaw66*r��Uvˑf"*�QK�C��4�[!Q&&��i#���	6�7g�ⵛ����
�Sd�Fӓ�f�sn��R5��Dh�VAG�$�[�!4}�Hi��.�l�m7:��	��,�uTq���F}�����t (M@����A������X���C{�f���!�S͵ƍ��IFq����i�&"|= �������^|��-}��8���/~�5mE�$( N��Ci�ԩS�`ĊN��3g��?�1�����{c=p"I�r^)�����Le���F�y�` ٍ�;<r���E�j�xM�q�b��V6�%r�D�������,	~�+�n����_8����@0�M��X�Q�{�0�F�n�YY50�m��Ʉ� �u��KUS�e�N0�T�D�92$y�<px��(�ݻGotCV~~V��5��i��	��wd�.lܴ��'6.@���K��H�;�����9MU3L]a (��O2hդ���o[s�ᔓ�E��3hj�PM�jD�څ{�� r6%�bAL��!kH����~ '����O�!Z'F�qt� %L��C��H&Xg�_\��|��Y�ع{'������8���,�*���4y�H<�_�ޠ��H��&!kQsu1?bq>��r
���I�
�[ʎZ8�?���ߚ]����G� �X,.�#������#��H�k�ٸ,"�����~�s���?�#h0z$gsR:�"33.̚B��Lx鑄#�J8�x�0��m��VCM�ڛ95t�8H9�����GL�u[���GL?�de���(X�S�ϯk:��k�3`����
�f�2"@D�����!b-&�ÏB"R%o��;j�YW���!�9H�ǠRV:i��7�ɤT��-8�!���.K�ТT\�\���^�Q���h��?,z1h���by}����|��%5:�H=�]����K�U�p�l�~P��עX�^������B�����8��ڿSy��]�@�;��^R�~�c21vM���oh
�B�$jل�fodi��mnv,~c�)����@�Ŏ�r�ԇ�ӆlN�	U��k��2!?���f�,`����3�?��_HK�Rk �c�1����@���ɦT��Һ����{��Nu�a]�k�3������Zfm�Q#�n�kv��x��f� 6�����ʡV�����''��aY@
�ϻ�mO}&hX��1.� ���"�>zCv�RgR��MP׾�y"�t E\�4ѓ>kt����P�B�*�0��k8F1#�c9��CîZ'&��]
��T���O8u�d"ٔm�QS%��ߵk1�H�����N>$'ﾛ�aϞ�E�rh�\�F
p�W^~U~��k23=-��vNW�w7j�&��yd�&S@m�(9v|��� �]�4�`@1���C��IY^W&��?cƞÈ8�{��u�Ѳ=� �R�� ggL���F!��{���֓�\�u�#"� x��	���\e�9�x�j�f<,��q"0���yzG�n&jR�ʑE=ILX,�U��L�M��6�ƶ����7F���	u�������H��m�;p��;�D��M��4SJGh�]O#��Z)�X|�4�J��Q*l��;��'��y�!�������["�����{�P��nD.��)'AQ�4�g��1��yc��b���`s��uc�V��fE\�������	?����b1	�&Lo=�ؚfx[�i�Jv��D��&���������QI�x_���!�;j��(�v��<����	YCD�h�֨�&L��#J%����*�i����*����ޑgBr�E���"{kDF�ȸ�H�Q=x� ��`h~��g��� v�&t��;`��ukL�]��� 7�C�P:��n��P�F-�����À�{����#-w�`*�Ӏ!ݱs''�^��Q#
$ ��YRCs��Y�&�S	����U�yێ���;#�y��P�A�b�f�_�N�l6�14rfϔn�5),��l;�bC)� lJ����âm�L����ؠ�7�ȾǮ`��p)?9ⱢM�;�R��`�Z[���gdd߰�w��%w�>�4�Ep"��mD.�����O׸0?'_������[dс�� ���ҘL��@T#~4҈���&�ϟ�{N�/�����&[��>)�.U	���!���FJ��4�$�����;0Į<yIƺ���;��r����;o�n�kެ�6\㈍
 �ݟF�|�h�&h�$1� _Y,.�1YQc�.G�V�[����=��I�v���$\�l
q*�lJ6�D�#u|Ц��1`x�i%Dm+��$�L�����z��pR��VQ�a�:K+���љtBgΘ�tR��Z�D5y7�VZ�3_*��tm �_w�:���lB �R�C�gPNi�����m �Q3ƥSit�{M*�5��lm�uf�#�Sj�T.nF�y5�أ@�xh�=pQ76$L!��9������,ǵx��q��kz%��F�}�7Fx�p\0�x8�+�fQ7S{���+�H�� *��&=��&����9�K7� ��
����9��#� �g��������ԁ�k]����5�[�3Z�>�(J
7�_aT��/�ky�чB�=[�8�h3(	/߁������K޺4./��ܺ|�i`t�4�:�����gn-I֭��Ɗ�բ<���_}���¦�?q�<��9��T���?�����o2��ix�niM���4�NkU����Al���]�Ig�/2�ǆaBñB�Sj>��4&��W��|	��<�}�bJub����V�{�&����O�*�Tr�k�[�v�c'8�1�Vk,����}�>��h�����c��ܹ��_��e�`m�4�0NLo�R	���z�H���5׉p�qI����m{�;N��Ƞ�dH�߸Nf-2��k���O ���3�]��,-�h��G���:ƌ�X�Q�3��]r��k����2I4�7��n���Z��N���_^Y1}�\������p��ɞ��Ѩ"�j�%��x�F��.���7�A��.�Ad���T3
>X�M�����C���`������`�:O��C�<ePT#p������
�jL�^�)o_�B�ا��kg�HW�v��'#}���C�I;l=p������E��:d��L�WW�L�*L5FM��3<��ل���2����������g�C�"sU@��X�6
�dFe����~,ݭ�=i�T>%�'A�C��n������c���~y����'�͌���>$�	ϨG��
�d�X#���*��$�Z*7�FOgXcv[EZ1�U���k:?k��*�xiW���a��raY�@*�U2�%�HҐ�	�D��ཨ��ȑ�b�+�Rmt���X���겱�kv��e��R�*��/����~�S!t�d�8��
��*#B��Q�����<G_#݄�����Q��ZN�2L��:�s�N.J��0<��9�usrwrf��"�����L�Q��T3KKl<ҁ��sX^���ִLOO��ﷳ�	C֊�Q&�k�x�g�Eҭ�;G��)�X[�а�qi���#�w�)3x���kš��j��+�-����:IH�흲8�&���1ԡa{N�D�Xil�$�-#z�h:����nF���4mYSo�!h`SL[���y��b���u��H\|��8�μ\�v�ĵ�.]�WG��Ů��E��մ��$A] "��^��>rZ}�1H|�ߑ�+��#b=8�jZ����?q�j	,OoP���2/���W����p���=�w��`�Ru M��P>�]�mr��n9{�u5�sL׺:�<o�N�6�iD1ۏ�)^��C�h��u�4�� ���Ls:TLK�Y��s���a�B��]dC
��W	"��P�$�=�٩q���Ԅ��9H�@M�I2�k�'���g}���ޭi�w0"�3,Sl��SLә`�:,��dmuQV���~vF���Eaj���@z[-G�2,3��4����ºx�y������F�hu}��v��ګt�0���b��70�	~��=��,4IPV�A2'm���  �>r�(
��"W~��:���z���];�]�r��7A���z�Z�{���|��U��\[8�s��{d�gt��5 c�G�}�sn�����C0Ea�Z#�u�L��a��/J0С��Kj�ܞ�%�fw�5x��ꢌ���F��Q�SAV����h�kϔ[z:��i�+�ޒ���G���k%3��L7a9�Vgg��_�+��7�I(	�QM̀�C)FA� ��cff�xXt��9yZ>�o�T�ȇ��./<S�х2S��	K�f[��m��dn~�?=-r�����O=)�OgC <���v�:���� ��g�uCA����?,��v�TU-�S�����jh�U�k�MĒ��"��m�e���zT+0�dQo8�~�:���A� }��^R��{e���|q�e_#�ڮ��a,����CF��{/�� =����\�"��ոY����d���=�3꣈��Z[����I�& "%\/ȊQ�
D�fh�Ȱʨ_"(@����_v��#;�\�l�n��x(Z�"N~�59�0h�xa(���:β�~cb0Mq����luQ�6��j�����H+ƚq��q7�]�?8s��k��ȗĘ�&���]]��\S|��l*���D+��1����LHѓW�^�:IՈ��8����������e A��4���W�<)U� �YX/ʍ�M4Z�%����zSF�&4:�HO���s[F�F=Hዥ*�W��/�ey�$Kk���iʟ1��!q�$���])��.:gۈ�����Z~��O�W_�ӧOɟ�ٿa$��}���s���L˵�W١3��*@|79;qE��ڔ�/��]�О�3kH�9Ri`��0G��Ԑ������.ޛ�9R��Y}~~��g��72B�4�}�\����5�h��رKy���0꩖
��ӥF2!S�����؇��O���I[r6�	�A��B��?Dص�ub���c�!20��5.�Çˉ�� ��f��.f���=k2�I����"4������.�9��޿�C��_lg�aD5CH�Z1�/���O�*0��_�H	}�ň�a�5BP�����Ec�;��Y�D�fi���2�s����<Nn6��+�R�g !@޿��Q�g����C���C
��뾣�9��mM�C�?�p��!#Pp���tey�O�5�L�4t]�$���\����T�t둪��$����F}#��P�dS�A֕o�bA�i�ow�	G�]��wu�����6s3"ecA7!C�TI�tHIo��Ĵ Z<�����	��L�ø9v[6*���S+g�1*Vc5����55��ԢF�KԀʴ I-z�5gӺ���m@��J�`m�ڱ~f�Eb���?��?��2��7n�b�&N/�Kk�8$����0y���V��ea�geF���G:!�]mM�`� �?'�5uܱG@��=(L�,�b��dD�x�	��t��(BO
l�_�����ϛ�FLB�חW��iЈy}eQ�/���^~��u3�2煫� 
����' �]{�"o�а:]�F �+K2>6�#j�ժ�I	�t�؉`�б���]Y]gZ���A��h{����I!�x��H
Le�Vgꍈ��FvI����b=����JQu@������t�����NiV��5�ǎ���^S��F�XZ�쏠9��ޗ`ZL���2��|Q�9B��c��A�����T������z��r��e5�u2��Y�
m���I��,��w?����f�d�A㘢�����C�j��Q�����@#j�-��TC^����S��@l�D�߼!�.�)0��9�j�YOevqZ\��"w��'���);�eztT�&e��u�Ah��KkĖ�w��1�����*�`�G�I����Ǜ�k�,*��Z⑥���Ԑ���y�M=�m�������o�yC�Y�<��c�j��C�42���9��˦Ԑd���_�a��[A ��J�bDyk��5�_/B�����t��gϫ]�cw���ebjJ��+G0���>R���ѽ'�����}H~��٨�.H�T���	 �V5R]�M~�=�ȗ��'�"�|�&�������psĆP
�-�K��@9�1ū9"�����瀆�O~�#YD��š�H�h7	���ɧ?�]x�������-� �l���^e�kM☶�VJ�����L7���sd
W�h8]�u��++`&�F"��� ��)�%q��jR�	�/�i��q����_�l���DD U����$�9;;��^�$߈�����5�j��3��Szm��WԐ6\�Kv�=?�7�����8���ss�L�̈�(���f�?ps�nH�%������k|nv������E�;�o���u�������_[H����Xj�&4��X[�թyy���pH:�daaP�gnɄ����m@�=����z�Kr{|JƧ8�&xrp�Cb��_������u��wn4JԐ�ݽS�����txxP=iY��u�#Ej����ƚ���	�d�u%v�ke־wUu��n�+	� 	�ARG��<vX��<��D̄v��3
�Ca�e��pxd;¤kQ�n !�4���wUu�[V���=罟��@QDmO>�X��Y�����]�=���+��r�Z c�2�S��ۢzx�E)�kO�H�� uZ�+�ZY�5�������A�~�7X��;{^�=J���1�����Q�)X�|�XDӞ��lkj���A��g>�Qy�Ǥ�/���(t	�on.��7^cgi5je��)�Fc��U*7�w U�jgw�_����g�Ї�2Fg�b:�)� �h�QR�P+ć ZdY��'���o��i1��������1d�V�Fu��"Jk��Y�ض�"��/��D���/R�HS�(K�����OK>G��1�xΆf1��q�4�I��5�.�7W�g�;#-=���Xʊ@��v��~�qvD?��/qs�{�rk��9��8C#0CGY��@�zU7���hF�������=���n���r��%�ė��P���56���7�*��d���uo�y:w�?S~��WGo-�Q���6Aʓyoc)�v+ІQ���ݰ��f2���\�JQN]�c5+�4̟P�H���e����/�h�o������t~]aG��9��@�O�g4_��U�椪P݌�u~�����k�3 ��Fk�����_�@
���& �p�oE?T333r���<R���C1���ζ)�7�j��$�#�vP_��H,-��V��1t"�1<<l4�s�e�ld�R����>YY��<�5�a�1��ExL7+�߇�흢v�vSӳ�����_�E��O��$�����/�C����ԯdw�
�uN���kV��)�mh��ƅ�6C6�R6n԰&5눒b�0���l�Z>��g�ȑ#�j���k�48��^׍�n���2�L&J
Y��|&O���~��j�i����d���x��e�ȑ�@�pPS>���U(�Ji*��g�|W�]��n ���*�
ho{|H��1�:���g|GD�`�JA�Q!&�`;���-� ���)�z�(��c�,������>ouUMGX
`[[�x@y�5��
^�>6fԎ+Ta���\+����z��̣a�,3��a��t(�w�w;D�^�y�1c�aj
��54I����\��X��y�Q/�'c
x��4R�iJ��h T$�n�ƚ��W���#�Íhʈ���|6����k_m�%�?*a��B��4���h��n�}���`�f��t�x�{�^�5G�*O�c�[ �C�/'�������~�yc��4� �V��##
�����~v�wVAh�)��h�~�<=:�۹Y�n�g�]PD����,,����^�5=.Д���hJ����k���|�����ct{<}欜?��@L����랎I �c�	��2����Hg���,gO��)=�x�i&$�~F������}�~`�uSa�I5���GO���韃�Rgu�*��)SON��ϡ� �R��*��D���X���k��o����0y�灆��y����x�8��t֍o��	�˵�0%������IB�\�KW������XJэ:Kr��\�]j����љI)co� a�B7WO�&�)(�J��
�MᆷkrJ&'vI�>���|������_�w�=���R��w������DZ[5� k��|�n� �9�{{�G
�f3<N��-���߻�é��r[��Q���,�s�V�M�1����drL�ы��	��� ���"#��J�8fH�RUP]˗di��E3:D�z1_ ��f��d�A@�'åX�7��MD;nӦ��6��4����H�`�mZ�I�) ��G|`A'Ag'�n%����6#��p�����R;7޴���M	��@�S��=�	��*��+e�t�wcx��z���9�3��Ce�EN���G K�Y��ҕ�7�ŗ���Y���\�(�����N�TJ]�k��r��ш?DxIA󷹉�~^�377/gϞa�u3�VOw���y6Ae�P�1�@���l�Z�<�F̿.�>��p�;STF����[�Һ%���Pc��z���?��p{ ��_��}&5
�d�D��2��6�]��%^_��cm��>��?���8���0��zk)��D?$�,�Vd�v,���|N��ϼ�~����s6�aް#�o��x!�� �@Ј'���V��������-�=��A��3���k;���(T��_� �xU�wZ���|(� �T+��4�-֨s��[(g���7��Q�[FP͓�w7��c�������c�֟�@� D� ��Y�a����P)��68�o�v�+�Z �H6%o�O�I �k~�TP ����h�2����cttL~�>G�&���d��<mu����PEU�5=�̴�����zF㽒ݩ���[����s�ʕKg����4z��N����8o�Σ 9 �O,��Λ�x��<}Y�7.��.��	#>"Vv/�QE�H�i�����'��ɳ2?�(��{��h�5Y�mZE��yըa�- �t$ܷ����<w|�"zA�)��}�lm�� �Yo�^O�g���֟�}Ĕ~N�$+�l�:}ܴ~nD��MS��y;�݇?�}|�~���zs잆��_ש�{��Cl��8H`��а�a���y��Y��zc~��X�h�pꕺ�.��ZPp�v�ٽ��0�0�M#��tNI���Q�[��nv�ձ���b�5�gGό����(.:�! ��S���ryN -a�aM��xpﶷ3�����{���& ǎE�=4U�׳֮�,ᘦ�� �����Bҧ���imu]~����3��������}���|C��:)L	�����ࠌ����=��8_z���ޖ�G�z�RFS�k��  �(�Go�:�5����u�v^��BQ�e�c'8PE�Uk:��?d���F�n  ҁ�^�d(���͸\�p�͇Z�q[���\��8xh�F-�3�3��}-7|��N�%D�	���vDx;����'���Mñ�#�"3�jtz�V���و��i���p36�o7�䶤����-_�6��z�e�^PD_6��ےDd�(�:�7�
~�{�� �<��g�DD��D�{q��E��l�:�0}W��$h3�F���~�G��2�E_�&����������2�߈5�M�����D2c�Z��	�M���+R�r�����m��e���/�V�O�dy��%	Fì� ���Q�\�w�i���	�0�H���얏=�$�q�F�XKe	M'4v@eB�T,�T��Xߘ���Dŷ����n��Y�L�aj��75Ն�sC,����_�6�~��겕YeT�:\4n{�y��h���6N4��!!������JH9딇����֐~ߗs���Y_���y���3��F5|�Y4���Ӯ��޷6L�8��s����kb�� 
Y��fK�=`���;��-�-���k���x��GK�� �R����%�d���r����qZ������R�]8��H��n�8�մi %�|V�D(!8��V���;Ucf��	�b���	s��yL+�pZ��u�n����{��'�+��_ ��?�z�o�o�q�kt|B"фg�Q�����ӽR�h��鹔p2zhu�:c��tn�U5١�%zel׬�4rk��Y��M u�Ґ�o%!�s��y޽@hxx�b���_X0�O��U�T(��3l���q�I��a���ش\�/�FY�!f���Έ�S���NWY�D�oL��ٸ��{� ���G���ՐXv�e�,�_����]���T��Ŝ���{'�nk�t����O�n�愿׍ǑW�0�w>@����W��q��l�3���q9��W�W[�41�8O�������S����s�05C�����[ln�>��~�j���r:����"���	嘞T�G��c�
��l�!z�G�O�`6<G7J�zCHy�Ꜻ0ږf�vo?hv4 �]�V���>Q��;��&x���Ԅ��| ʘT#������'�d/���䩳m�5��JÑ�����xF)�mg
�p"�LmC%'Ǎ�l���]	F�RV@F�2=�_��A���ZU����F�[r��#LyS4�k_g (Rk�?Q^`M��L��)����9oD�� :�E�95�0�zL��h� {U[K�|G��I������"�2kzS��
EB��d�� 4��"R\v��k2�{YYZ�M � @�E��Wgj���u ǭ�Z{�w:nKJZ�V�w�-C<cW��~�J+65�F���yL>�]`4�i ϔ5S���cG��:N�N�<�wz~�L���n��^��-S6r�9�}�VG��j#�W�07J[���ϻnR��o��Q�VeT���`1q�� mʍ�������kN�|�:Ҫ�9^�Vj��שH��9*��Gq��oə���K��7��"���i���,-J)�!�@�*���ݚ�D{�P�����n*�5N��ĴL���t�ԙ�
�s�ҋ/�Z��?�	9y�|��_��/������p|�T�о�{97ߤeKS�����ģ�ǂb�6|��P�eɄ��f�����njʳ��F&�Ge �=��fw��B$�Ͼc&�t�"�N����"���q:���-&m�t7}�x��u��Y禍?y)���Q�95�vv�w�8jê��l�����������k��ns+ښ�R�ӂ��l�;��?-���u��mѹI���9ކ-�y��[G�Y������m��h��ps�D�۩��-�\��3���[�F�Us�Ӥ�!�ptk-to�%Vcȱ����V
��.|`|�7��ػ�����}��AOO�r��p�ޥ�z����G�	G�2�kZ.�OH�5�O��4�>�� C��*H�4�.�-���e�dK�9�y#Duw*f6�ꅳLM{�Ҧ��XZ��+ Q4ݖ�Wes;Ka�{����~�]L'&'e������<uJ�F����K��o��j��� MQ8���c6�z32	s$���3��(�#��׹$N�%c���ֲU1���"�Y~ѸͪA��!�	57p+��N ���Y��
�D��*���k赍R5��b}�9��rf���ؿ庭�r;@�o��-�!�훓��	�o�N�L��9.ݾ�nm��}�O*�ubyǽ��Ag&�~,Sni�P*��A�a`�~L�ѷ�=���3�[���7��{��o)�`w�6?�#JV�`KS�^żGn�7Z�G�41��NEt6��#v�h��v���4������K?V�ې��Y:f�?p�㌋�cI�{�!�1x�s�o�e`pLC����lE*nTz5fk.٤ဆ#�Ser6(++k��U�L�
'��(��Q����c������榬��R^AC
��:@}��0g�F~u`v�1�@w�I�tiTȎиGSml(.��i@X���5�ё�x9�Qk���[q�^$�Ov"���a��u�k�,�!)���9C\�)�5���&W�\�hz���AnX�ԤD���~H���:"N��������x޷~��o�i�s��ρ�|Z�i3��A4yC������3{��h������Hkh���������mz�t��i#gk,���u-���40�P��כL�A�GD
�s!��س��������_��BB��d���p�t-�u�| ����I%S28:)��xH�er�:�\�,8qx�� ���#�h$Fj�O�xM�%�qP�M����g��,Ӧ9�:���g�^��a��j��R]��٢���@�Ś��n&P%�z~�(Ug;&���%~`��4�INk��ڌ�*���@�O�l�<P��^atL�68���㚨�/�p�&=�VVnʱcGdjj�χ�>������C����Q����~w�ܫ��r�A"2P8tZ��+����s�R��ކ��F�n �m��G~h��<����5��[_��RV��6��"��H��Z���\r��y1���E��iвl�j	J��C�.��o�o�@� I��s���G�xRA,I=�'O���Aj��P�\�|E������L�H�V|A_�A}}������0r�k�E親�1�(�Sx ��xmG6׶%���Fɾ��Q�O#�:�u��.��Q�<GV�N���z?�0}����)R��	w�u6�`�U �k�BÆ\��h8��viqA:���9��ʌ�#��=�ʹ��^��s������A4�F�]\�VS[Q�m?�Ѧ0k�F�G8�c,h6�v�o�3Hiu-;����[�9��y��A�(��%����,��`J�����G?�.>�	㎈D�V�Ƙ���Z�0�����.���7�{��)=|'�����~�W^����_FG���+��������=YX�!��?���D� �4 >"Q�2@��{�����Pc,a4S�9��eΊ����Q�neyA�r��=���$NH,��6@�T)p��V7��&��V���j>y]S\7�)�X(�Sʯ\�Q�\5��W�A)ēs�9��g>���l,-�����7?�NI���X�^����덐�qp���uK���#� ʵT�V����W�g�rc��ب���S5ݹ-m������E���ƀQ$�k:n(d�@l�O���X?П�4)Ӑ���J7>��H�<��_�,޼!G������?��	���@����r���W��瞧�@'ʫ��O>E}�^�T"!��KuN����#�s�q��֛����9�zť=�r�-ٻgJ���G��C����8��u���� ��|�6�M�z����_]�0�V{��!y�����Ņy�nlmlҾ`;2:&�}�3��E:�g�<��c[Ay/67wÈ�X;�nj�]w���T�w C�C�C���'����[�ݭ���-y5T���x�c0�ڐ��y����5:��[z����DV��ћ7��K�r���2<أQ�(=0�5^��� �쟽^��֫�����Y�|�!y��C�l�JA]������?)ܿ��f�X �J	��r�����_b��)'�PI�k�!j�(���_�u�G���9�\�zU�W5�P`�'��WOHoD���_��}��җH��F%����sWds{Ma�ĒQ�f�b,��v�>`G�&�Q�7)�vdyq^�ɸ�kԍ�����zsNv���:Y@';�}��{��ö���������v0��!��;��1��)�$|����X�`�@��E3�9;&�l$��ΰ'��a��񵞩����֭ ����?3�cF�"��5��z�s��k���g�$�詄t7�.ig�=�2LW�M}��Y9u򨦫iy��$qF���,?|�E9x��|EA�GY�W~��\�zQ��C�=|�T ZY]��t���9�B<o�g:�ѨU�'������׏�F:ԿW�F�%��>x�!y��dblL�Ţے\<wE���Kr��	�i4�L����R��T�6�����j��8��	��3|_4��]��yh��
%*c���	��z��Y�<�{���u7,;,��uLD)���0~�#B��s�7Y�k��e^�H�N��#�`��M�(Ց���AF���A��7�����A�Ԥ�����פ[)O�1rm�������-U��+�='�<,�¶����7�X��Bޤ�O�\��ET�  *G�����7�l=��k�e}cY����d��[����7�/��Gr�FV*�:g��۔��W���9�ٳ�t���rs�,������@�W��Bt+�R4��L�b�g�!�;��"��\���ݒN�eS��Q�p�ir|\R	� �X�/y�Z�GyT�GGd3�e&5z��mQFڍ�XP�)f��"��C�L�a�t���9r_�x�i�'S���g<ˣd?���
`���{_�9��8q� �]w�rm����n��N���ѣm��?<eD�q"�0U��t� ��ψ����P6�jҨ��f7O���)��ZN���yY7è~�4i�%vԴQ�q��Qh�|[��v��2.�E�u��KK��nIT���U�iTF�,rt
,=�RU ���Jue��g�e��*y �Jmnɮɔ�{�}�E�@P*����Hz��|�=7�Q�r3$Y�^�d6�������_|_f���\��O  �cD�P��'�J�!�n7:�z�����1�i�^�g$��t**�/^���e�wH�N�
SS�Ӳ{vVϻB:����|��`k��mvx�B��M1�
�Y|�J��-SC`7���	*�Ch� Pl� f���fjږ�����":�Qö[#�`9���5؁{Zā��[Ų�M������Cکjj��?��*
ULU���F��֍ E4Z	jtAr
�>a��	��<�j��٢Cv���%��0�\3��@3�֐FzcT��SQ��ޤ�����b�0飂����lN��,�4�]S�u8E��ݣaGvH�자��7e����Lht��nA<�S-h��ய���� �B8]$&2�	 ;��)�쎄`Ά��^�P<&�#
�=lH�A�O7���	�ru^���*ٝ���Ё�Z�4���	���lpZ([�\n�[E3ɸ�6dm#'��;Tf��I���P"{ϖ�[и"�
����g"}M��@��n����]�΢��e��l��>+Qc�:�MH�X+���(4��+�UŇά>>�h4���jce�����Y�#E7�jE;�_�RzP��-nRM=1?=�p����~�׺'b;u��j*䫬�ժa:����������F�� ��H/�y)�Ϻ "��F�ui�˒�m�tα~�ZQ�[+��pUy@�SA2��n*�̶� s�4��w+��oK ���а�&��W��!ʮ�����R)�U a�d� �L5��k��#��@7��ܖ���Db)9��Q�z�n~�/A���(�d��Z��Z�hp[0�YlF0�C��Yc��.\#� 6"C�����(,s]�ՠJ�6Ƈ_9,�cC�_����L��Q��@����VSw�%�s�֥t��G�,���5�f ��{E�
��zY"4�T�H���tZz�f����3���?��C�L&'�lQ��z�G��1:EDZ���tHUj5�DZ�SmU�4$4e ��p����k��vh��$�c���<<�"D�ґFN��@ j��Bj'#W.]�`6	`B8�HV��z5/O=�������G���G�P1�T� j�eJ�a#0V�E2�;���������iD�s8�(1�����dlG��ʊnl�*Ĕ J�s&{[z�J�5�*I	 皡����4�l>�,�����Y�h� �8&�/�ES��N�il4*U3�,n�
Z1}��9s��^8?�Ihާd8o�������զo�4[�,��H����� �i�JuU%���`2%S�C2��kY+e���eH�a �W]�L�^B��@RrEXשQ�* T��� �4�X�x����Ի�p#�5Z��Ԡr{MS�c=&���"������FA�Vc65KW�7�22kj\u�j�7m����K�|sY�웡��s���D�������?C����M�4|T��G����y����c����#��oe�T(��
++ƺ��S"]*H�B��ry
��`3ri2�o* �i����:&�PW-�:P4۔=�i�����tGӚ�a� M$�:��t"�>I��h=�_�]��nc��#ac	}��Jrn������?U�ٷ����h��]��2���0"�MX'�;�n�"����M)4��7$��d������~	5�o�����aI��F30��C1��Qo��Fu5�@��������TK5�`��P���B�/�g=�"n'�5SW,��X�	�(���0#]Y�!���7��(ć�;Iq+�)� 4�&��aU)o�O�o��O������)��]���3ҫ����>-��{T����k%��r��)��W�Ϩ�FN��eu;'~���Z��t�9	�&S��4�L��PƇ�|O�H��JakRӍ]}
�*Xc�W*k�m�H!�u���,%`��7,�xd�Eҵ����P; ǆ��(&���>5=�*�F}>+�֨�X��Z�9&
G��(���*�<��n����������]|�]ZH���q�mP��y�����=6 ��I	ꍔ][���2%��F7y"�Oid�nXJ��Ӳ������(vJL����5M[K,��13�԰6 A�-�=ɕ��c�`��m�Y�\[��w�4,D��ͦa hD��Knsθ�j8�ZގF�hnA������_6��R��\��S�L'�`oRPd}ÕW�.ǎ��O<�1��=��U�!�;�[f4b?������ʚ#�����X�8v�+	I�')�dT#ㆦ�e���o�'!�����v���V��U�\�t�J6��h1�RA��o�r��؋�㲃o?P�;>���"2�L�	��C!����e�|M�+�L� �U(���R2�����F��v������*��H=��;�Z)�v�PYj��eb�O��R/�HF��:���R�OS�b��׬J�X!��C~	�1�\�-��Ԅ�ECV6v$��+�D}jN^*�Uo�h$ҲG����g�����\���E����Ay�C�PBj��E��t�CA�=�i��&��ֶ�LT%=���M�B%��9��o|O{�1I�&�²���k����\�� �d����i�F��F�u9vR�n\��tXҽ�g�RG(��Pe�!q}}�)��h��$���jy��v6W��P���B�o�_��v <���5�{�����rT��Z�0�pZ�Zd���3L_�0��=�s�j|�h���Sئ�Z����F; ��3cù$-/�:�����hw�5���l��tߝZF�T?�5t�1ڈ���)5I%�2>�'��Ov�W���Q��U�H�֊=��sUS�J���˧Z*= ��A\�V/����hWV74,h$��F�%��X>c���&�P�Q��w�X�P($�����;��/|Z������C%0��b�K�@&�g�%�
h�Tj*� ��i��8�(�������IE7�?������|S�F�i���)�/\LA��˫G�3�K�%�I6�(ۛ��ɞ��dO�Up^`&8v�+65\�= ~ms]b`�1�nn���w���yIBH$�
<��(��wZSa�2�i\�(j����uQ��c��v��3�6�>�x4��1 �D�Z��RWS�
��z�_$~\?L>�sy}�6�j�2�82ܭ�v�]����Z�О"��N,+�l.\�4�7M:���@����C6mbt��sFA�iE @p4b�f��e�@(&3�&�Y^��L��)MiQ_�폶 Q�!��w�3�w��P:TV*�[�\*�W^vM�ɣ= �SC�%�΃�Tm��B� w$�n�	p�I7L �:�@�\^ؖ�r���y�M	�Cu�"����
(�v�|�kg�_.l�e��7�W�K���o鵰J	
-�e
��i�p6���/��9�b������H>���}��D����ս�`��E5��0�xL���ƴݵM-�U1�>�Gx�y��\a�gRz�׎�R0�`� l4��~�����Hu�T5��
��2��-��?�ewt��	�̪�?�j7�|m	��zci�״q���hz��Iƒ2�pS��㦌ţt�lj�Ҵ��3uP��0�K��L���c262,����k����p`��1\�r�4����ԫ5F��'�e���섌P<��Q�f&+�[[��R"���5�.H� �c����Bg1W���+�oJ4�t_��H,a���ʊ�ޙ�F�%
��O)��\DVW��v��M	W���͢X�ج�b|C�z~���>�ѯ�<$���D��e6��A������ׇ�Є�l�F��O퀄i���ȱ������Q�E��������o}�`�pD�(}@t|׺��H�֍k�/!Ο��^��3�zjX�'�;��]w��23� ����u��&�"���F�9�)�po�$�UY�Vehl@&&&dee]ַ3��%K�AD
���A��������$[���}��5˥l�pLm��hݒ�k�R|@��c�*�79@�&����zD~�ҋr��%SkW�z�
�x�d2e�,(e�7�2}��)i�C2��K#7�>�y`@W���=f�S�4��b`a0=(�ܪ���+c����hna��Z
{@�T�ОD��r0�L�d��������+��s����aYdyy��KH�1���R=%��m9#����By�� ��Z]|�\�ݴ���j����HU�!2*�z�)�f�[�
|�t)TG�i���]��r-��Nw�^>���
7Կ�(�${$��m�)/fc+#eM�.�L�lhE�����H@#� �/PjJl�D�i�n�#}���1���$嘱F�fH�����c3�M�(Q����-�QC\\Z���e9w�<�"R��d�(@�X,�a��IIY#��Y]Z�"#���P_Zjn�)n��K4��R�mM���<� �k��2�o{D�|�K���^���ߔͭmI�k�잕���Gz��]P�^�,����'�3���������~�i����X�I���,��`��IX�4���
�o�S�ƨ�m��H��x3l�5YS`.6tC
3��\�nc���k�f��%��\�DI�:u�\�t�#�}p�� ]dV�P������}��'���Q�VD��$��0C�'K��T�@b�
F�^*i�F3(�w��4�F�4͵�{t�!���%ڂDz�ͅ�X�sG��j��R��&c�١��h�s:	7u_o��XN?.5�_��������E>Q��������)x^�r]�|㨜8v���H��椡Ǐ2��FqkaV � �5���l��B^t{t��FQ��-����G���ԙ���r��ٳo�<��c2�g��ټL�O��ں����w��_���-_6�!�9q�F�A�D��^�C�Ï<(O=��)��8�Q�}��������Ƣk���c��zK��Вڮ� �_�v]���dgv)�XzHЧ��^�H�D�'�H�3�CI����2>:(��2;+�,����i�;�Ծ���m���'�=�&���]�D�!�j��f4�֔�ѿ�#~v��FH���M;�	^cP�5����T_�vu��	�=&���Ǻ�m,Ɠ&�S#%F�t��t*��P����e�<����X�qM7W�{Lm���2>1!q��NNʈV�A=ߢeTz�R+oHU�uvz��{������+`zR�_�,/|�{2sQ7����so\V礜J�@�_{�	9��^�53C1keM�+M�����]�����}G�)�"���� M'Y��33)_��/����$S1�_��7�x]�� �zAv2[���J�Xoo��1�t��Y�8���M�GpP�=��T0�<���q�r�Q{�VaZpE�
���N骾ޡ���G�]��z\=2�י*<S��f��u7,o;Pa�]:4���l�]Z�Q�&U4���_)��q�p"%YM��w�"�t�]:�4��p�֛��y6	���݄8��/��&-HE#�M0t��qM�뚎�(�a��|�K���^ j(>~3V	�w�JhzI���
Ԛo������y�M���i��I��T��&����=�я|T�I�v���#>��ɥK���BX�н%��Ȑ�����ߕ��y���T@��ï�F�lDt��=��>N
ŬTA�*UdaaIy�P�F�ԇfW����k��(�;(Z(<t�${�l��]r��Y
H�2�*e~n�b!��tP��-� ��I��(�����~�-@�G���Ͳ<�r���y�IA˔����%I��b#<x�=�ӌ����(1�[�c��<��hw��-dZn�w;i
�X�Q?o�:�c�b�\N�5�����q�|zIjSf&f4��IA����޹AO�u�<E,0:��얂p�@�J�����|��FY��*jZ���y�3N�H%ۖ��L�GXbI�^�Ԟ&y��t������ge||L�}20<,�Tʒ�CT��8�����%W�A�I��/��CT��IF)=1�/W/���_��F ]�ɧ�k�(�|Y��^����������{S��_���'>�	y��4�����m���&�^�.(�wӾ�݌��`1��zsP	SK�*B��T6[��^��vV��nwO�ȶ�����t*E����;���p8!5)<�� ;h�����N���x<�+6�r�<�"h���z<x��<..���B�ܘ��������)��ƣ)xG_��1�TЀ����h����!�C	Ih�ӃA䂺#��Q
+V�L��*�1A=ԑ��gV$S(덦)|	b".m��
$�XX_�B�"��9��������Ŋ���?�Y�0��_���������S��kRz5�p"M��  G���A���sB��������ʎ(���3����5�t�~�Ԓ��a�c��cÒ�ղ2,�+�� b�v��	���`�lnmRhv}s���)]:|NDވf��Ɨu#z��19~�^�!Iă��������db|Tz�)C�g��y��o�)%t)q��.�F꣇��!  �pIDAT���)���!�wt|Z7�4G=� ,@ӿ,J�{�4�uS��eS�T��o)�///S�,蚲t z6O��;"�]w�B���;I{�V+�Ǎ��m�#Z�K2��,�������8VV�5���@Ta���ڬ�Abw4�O�L����9�	�N&��lLW��=��6rؘ����[ �V�3��xb ��Ύ|������z媌��?� �t�	����ɇ�5�Chڠ>X�sASjeu[ʕ����J���������`8h��~�}�A�U��7��h;�r����U��YwN#{l3�����1��e���Sz�k��Z�!��Z�o~�*C��{��i�����1���Վ��`����3���WŎ��eY��:qꂂu���*s�R�e�?�&۬j�!zܛ�[%�����^%������LLNP��z�j*3�]�uw,J�;<c�[���4RA���ݴ��-�!�����)M����.�+Wd|7u��<uꌊ� GYoʼF����䋒-�P])�r}aI��/=�=���I�V����
N��q���Rls�W��W=(���"UnѨ�AFZ�� ��y�� �`tl���u���A����G��%F*C����6���1��&��ڸ\)1��ݽG�roި�6ꦋH��D�8�c�=��d("W��ɿ����|V4���#��9uT�H،�>]́�7���i1�Y�X[_�S�N�+�����i��˞N*Fk��sO�C�Cbqi��]S266�H/�@��t�5��{���G������"���h\A� 7V��&���P���S/Vdce�M4T�Ɉ����-(���L}&WP �h�|���:iR���FTS�:����c���2�t��_��iZO(?��Vv�<�?H:RR��W._���={M�
MA3^B9B#,4R�0�L�%=�^�'J�q7�#�������H�ߔ@�@��㬑S
n+�hЬhӁ�A�/:::&�|���7��ݠ��ˮ�D���m�/ML���i:>� �C�����%�ݦ�e�zBĈho�p�����IAg����>J�o����fj.��۬��o"e�)(�FtS�B�VVn�1�q��ôopYE����u�,hF��@�:)n(tx��`ZT Y��I�rE�oX�*�z@��ÒY[���Vn� �U �1�y^��H������[%mgKO���� Q_�f4����D� ͍�>J��[;d@4��Ev�''w)X��t��=�l��	 �sT�!R��@`Ѭ>�33��� ?�����`�u�t:M�h��}�ssr��Y����R�H���$�7(��#�?��S����/�B'���4��<���ɢ�I�:}[j��edl�Ǉ����ȔО�oĜ��L�����}֫���[�c	����R.A����T�j4�D <�~i�
Szd���>}����Y@��@AS|��B�ګ�vWw��}��@���#&!M 4&��՜ =�3���\��lE�o|�}�78.���4�Fs�R��W�Z�h�@��P��eQ�7�RD�"�����@��ƴ�\�5��H=��� .�%޳w�؈� ���l(\c��	�x"����(W�^S��򹦧���g5����y\#�=T;*�)�8,ԗ@����\H�<�	�����:mJ����\��dx�.��͵`�S ��\u�=/G7��lP�LtQ!]w}T��!?��*4D�FA��[H}~s��gOM+m�w�֙	��{8vxc�����X()�\��8[��(�+��F�x{ �Ԙ�
�t�]�L�.�^�H��dD2�$��G���TE��`\V3Y�9zF��22=:*}z�j:�38&�UpAmΩ+x������\��L�㤎�r"�&Ђ��H��r��e�I�G�l�kŝ�#�L�[DoO���vϻ�5>pŬ�S� 	�ǎ����v�@?�+ј�4,<WAA0�@w��5F_�7p�hѨ�F��C����9ų��$Ǐ�" nnlS:0��ZL���s� ���ceyEA�,�w�8�
&���\�~��EQ��!�=�9M��$�}zm������4��3�"�L���P@�8sF�M������Í�ؾkZ�\5+-��kE�+�:�Kkuh�!sP�R�Hn���7n�����1�hQo-�|���%swu����f�6���O޲#�d�ꍝa�'	zn@��$T�k��IK�P��K�r���@�р$aq+�"oh4��¤���4� �]��0(>~���z8��T|���f��Z�&��Ws��~�~�F4	N)��f��FFƬ��+7oޔ?��?e�z�=�ȃ>$����Jjĺ� ���7����_���.����'����B�A�<�'�7&'g8�u��E�� 엏}�Y�^�xAR�^I$���k�sG�=�G<����!��G?*'N��4O;J~?f=tGs���T���~'�4 �<7>���*F�Yl�! z�:�ʗ_7���1���f��Q���G
�R)�34����Wr��d��cr��1Cء��_���]��r=�s�l����6=Ih��33�wq��V�F���ƛ�in1���H�Rk�d�\�B�[�4�.�<�H�z=�`Lo�@�L ��A4�g]J����\��F��=��N[$�n�~���Łx2$����n���%��S
vQy�ǯ8����إi;  �/�}Xy�1���f�v�&Z�!O�ƂY|��� �Y�p�~��tzP_GS�`TN�8%�O�����=(�����%�O#dLa�����w�'�u���R t����{����r��
RE�P��>s����Y��O���y����){�;6����$��? P[6$�˒�O߫X,l~f��ⱨ���u�G�.��p������������*��i�jӟ\#�F��flڬiR�&�ܠ�H155�2���Ѫ��N�D"����B�iA����A��9���(:(�9�J�����I�	��Fk����X$@&�rb�?�c
g������˿�K255�T�;/� G��)�:$�{f%�Jɾ}���T��nʵ�E�&�I��]�S
`A�-�a;\.Kf{S.�?'�cS�NB�0����QtT�L�Uo�O�Ҥ,..��sI��&�y{���r��%�(<���k���#S$5K��3A�- 4�w��Z��U�JW�ϔB��J:Z��5;������M]���Iy���n���Lb=�HA����M*NwY�\*����a.�^��v�]�0��^��Z�|�e�V[rm����F�u��Ԡ`/�7D>!X��b���
�6�48-���>1R?ȼ�l�������p#Մ\��r<��{�=�S�' rC�
s9�0����?/����������&'&�z��#3�>�L�#G��_���
��<�$WV�u��I��y���%�7oR�	ͥ�F>����E���x$D�d����E6�֩ݹ�����˗/�9�;��STP���W������*�\!���R*�b��h�Z-�M�:=�b��
E���c� `�S�^[��(Y�GAqg����Xq�������Y2��b�ANlOO�MCqK�wG�����$��-��>$�*؍G��X�6�{�:��g��.���N5�Ń]1�v	�zyp3!t!nLȲ��u�Ψ��1,C(1(P�T&(�#�5Fnm������F��}~��5���=��g�}V�?N�9L�����+�s��B=UM�	I$��
����cM헾�Y)A�T��K�rce[N�8)��_���D�0X5�մ�\�I�Ff��ϟ;��&As;4��mSl"�7��ob�����U����Ή����6���.j�]eT��M�Yf��Ш�R��T����azL]�cCrHCjқɸ���$�
�W)�� 0����|hBUh�\-V�G0��u#Z�aGΜ>)W._���f���W�V�Bѷ�۵﮻`�-���
�@�)�!�S~��6�M�)�۴4�I���eF2!Mik0|��M�#��NTc�LxS�2����c�m�fc��E�^������G]ӳ[�z�7T�p�����^8�z+x�x��̶d�y�d1�� 97"��)q"q�h丶��x,!��q����U�(�qZ��ʚ���d`hPr;�n�{p���INS�K�.�t'@�op`��hd�w�,U���@��^+��걆}l� �2�5���2� �T�)T������0�r��tp���qqZrb��uۊZx?1������oR� =oB���(�/��_S(Д��m�l?� j~�-8ݮ}w��=,3Y�;C)r�>#m654�P�Ff�ҍ���>�t Hܬ���h�5]4�� ��5Q�aM��Hoh�4�na-�����!|�n^�Ȗ�;�H��gzf����[n�4��`	$<���*�}��(7�+��ܜ��w~$?x����R⮎h:��}�2�kV�5ş�zM�
R�j���EPֶvdG��������o�������EAQo�֏�ED���)�+K266"#c�4��Ea�Q3�Z��,q�itd@���e�4�a�:���,�����*���b(uc�t�#��M�5�j������r��A!�Ƅe��qI&{荅M�o�4>�ʲ����d���,mLÏK߻�gNq�^�;k�]wϢ��{��ԟH��94[�EM����k��ҭ5,-H(�'��`AiBD��UܘM�m�k�	�P�)-�R�#|�9����i}>_��5�̸"�H��ЪT�f���|"m��D1�'����ĭ�'���QM�ȞK���EI��x+�d�9	�c�ֈq:�T_�,\�*��M	k*��Ge��eN7}�gE�rӾ���o��m{ �ߣ�!����8��X��v�[�R(DWXs���<'�~��gvFS�$M�t;`� �&ۙ,�.���f���,B�TP:@��M5�.0�߿����^ш���7<4,�v�"µD<�����oȧ>�I��g�{]�n��da!�pM��]��~���{�lDJ8I��Hj$%������F�e���ڍ�ih��-���J h/b.ф��~#����D�do,]�� r9�
�;ۮ���, �b��itԤ�MSzp�V6Ro�����Wސ�g.k���/[�bz*�G���n=�̓<�~^��%���f��p�8���]Z���uzTM��qh*�>�67����Ç5�+�I-�:�S���`U����h��~�҅˲��,W�]�a�B���3�g��CfM��q��:`C��`/��q�,�$�#z�	�I��	�W����3�򑧟�e �!��^�����oh����Ul*E��O}S�VW���ƩϤ�ٝ�n:iG�R���Vɫ����.o�Y�!�[���[�[�u��_z��1�����]3�IKU�e���E.p;h�����r쏚�� TѬ���&��Ss��mnn���yE������s�dD#)�f�}���f�Z ϋ�F(����%KR���ɓ�?<,�����1���3��(i��\!'gΝ�A]*���I��Ȱ�s�2 vr
��*���=�N*�(w(�Bp�F�c�}l@���o�1�_�%�җEx�~����_���(`��IngKN�>F��i����U�p��d�4�������̑��`�( ����?��n���*�ŀ�/x[!�����5Y�_hm�>]�~M�4
ǘ���"�z�A�цk���Ҕn���޿�t��=k6�:���F/h$ Mk�����B|t�V���ռ�z��=I��o�P\K�n�a� � &�:]���|���z�~_[�pZO��ɱ��w��_�+)d�iuܾ��ڦ�;N>Λ��4��H0ɆRVS�F�_&>&���g �Kpi:��YPPA����&���b&#ッ2�ꑓ��|������f���X����G��!�� i�
'Ht�j�����o��&?�#�X�����o˸b2��i't����U8�f6�7��v����10;��#��xWW�4r�SS��nc�6"=ɔ8�Y>��j4<&�|�V.�h�Ʉ���Ҫ$�f��a����3u��3��J��X�q��B ,u5ի��AҕH��ޥ&{L�ʦG��ZR>c�k�l8yÞ-��J��1�aRM��G��|A~�N����)�

��&DJ����K]�����j0�m:������h4�W�M�)�dcuK�#)��,�B=�ڨQ�/�쥈G�w@At[��R(U%�9/gO�.�ʶ^X��O�4���\�	꺜�r̄��_�����s�����������dht��=P�@�������?���>�Ԩ<��1@��ѷ*��KS��5�rbJ���^ǊF�
�
�v��f?&�>��ǹ�5I�rS�}z��%9��+,q�)Ծ���7�A<�8I�U���Vˎ�Q`���>[-�Dn�D�(!fҰ<R��u��&�<u� �):��ڙ#�cPף?:)P���X0��'ma���������_��<��}�yO6"$�W�|�Ι�rټ�(��˽��-G/�șk���G�iJ^A��Ɖ�rr�A�.�~��zR}�g�q�xo\�,3������}Q;v�Mz���⥆�Q�
T�<��_A��[M���Kr��%y��cK\�}!�tmQ�rU��ӟ���Iq52�"Wv{C�6��2�#�Z��W�H��� 
��;�7
�
���)� Ʉ�ĵ2T�,H��eH�ZP���)	h�|D�>�᧸�A�5�,�8��B�FSw�5˔O��f���\jpb$��
��9Y�%�KɥMKj�0Z���#C[�����;���B�Ȫ�#z�B-�;�%H�Hk|b�Fl�������/ˁ�S��i�kK
�ث۴��օ���)`�������/(��s?E8k�1�4ڍG"�H�"��,
���]����������K��	�j�|�+k�兛��0nڪ/��f��є��a������_���+�}����Ï�x����]�퍆9rF^��r��%�4�r��y?E��
��h�1]�]B���ֻ&~#VE�~Y�pS�H�q]���ln�8���ݻ[>���[Р���8ͅ!d�]B~w��}/�O�5b���!΋���r�Xɵ��q7��6�:K�f����z���SǀPH�V � ��o0&�VjR׈u��~�M�jq�������}���/{ �;���ڕQ�B=SR��+�SnT�RS`GQ���rN#;;�^q�z>�)X$�u��� v]IR#5��.�xP��i$-!�<k�6k��,ܔ���v�0ugѴ����src������8y�ͤt�_����Ѯ|nG��Vem���샜 ۶b$eڟ$��m/��� �'D��w���8�a��㗢��A�rŨNa V�P~�KU����ɵ���۳[���_��}�r��e�e�c5���"iw���Խ�HE�Y�~e  
���z�ۊ2;�`��޵1�k�l<m:���[�j���=���r�6�(�&b#J;a}�R��9]�E#dtt��(6��e��_�z�fL�v��Bs�-/����8e��"��й�x��܊��,�ԫ�8媔�y��"�A2"A� �\�Qdg{E�}U��П���0��PJ ��j�����>ޡ�2����I��{P�G'eyu����_�\_f����@8$�T`�5�n�7ȴ TÂ?�U*֊:H�D�4���&
 E���P�yx=9��J��;Q��ƣ"��&vM��C�����-)+z���s��YQ#"�8�ɦ�+�8�Z�wp�x�$ ������jS	� �u��(�iB����:��}M?����m�y�j��yp�#n�J���C�\*�f���>�P}G����7Hq�2�E�����_�HmmB�= 1�"�A? 2�-��~U���ŝ�8
�9�}{�QR��_�j}0��;��F�er� +X	�r��0�P��W��J2"�ajj��ciaN�w�<rh��.]�����^�_�,K��$Е��*D_XʀM�/����=�H�ڨ��_��/��`��u���n�$�dȗ��s8�)y=.����iT���{,�3�s����GאE(��a�7���3�z����/�(jȜ�����6|�P*���.��'ehh\S��zݒd������m�[wu�{��NB��>~6½�h�'�{)n��
��`G�i�<�a8��ƫ�G�L#˹�Ԋ5R}0m�)8@�q�"GA����3���O6m�
:N�˼n���n���;!n�XC4��D����}M�t[~������YZ^bC��}��/�|�Y��ѣ�da�&��N�>#Ǐ�`�(���`-�9�$��Py
JO(&�[��Xa';�Q���Q�'$��p�������,/-�~82<B9=x��-`s+C��/Qe||T��<����4�c��ݑl
�Ak]]�/U�Ɓ�傏<ԟ(`b�U�|�L$�Q�x͎���F�h��sA��I�D�͵�*~@�<S�v�
��,T�K�ۛ��#�I�ƽ,U+� ��2�Khg����j݆������e��Qp��:�	E#��$��
�bV*�-�L�sk@0��ik�O!'��g���g-@?G�4

i������o�Kb�S G4Fܐ��I� 8�� B'9��J:WPv(Sw��i��y��dxhH�^�*�[[�n�D?5�i����Fɳč?66.�}�r��YY^  �������p�Ǔ�k������`��o��<��C���"�RVz�Q�=�K���#K7o����{�g�wry��ťU���D�v��� �bL�ٸ��[.�9%��P4k��;�����ۀ�<��o1ց��?Ry4��E �|��
��� �׍�x4�@3�J�z+��%:��X���!���[6u0��Vj�N.C��A�uܘ�*�Ɔ���Z-d�Yʳ��%�QU�"=	D�f��
\��
4~+Z;�ހ�P��C�6>�����(�'-��&��4e �� �<�*�H�$��������dOJ�VW���s���dttD�FGep`���?@̀T��_�홝��~�323=������lmnH��;x��N���NHO�G6��ׯ]��=��:2����v횐H((3�vYF���4Z�_����r��)�*��Q'u|�����Q�J�`�!�DKz.���߂���j����@I�w��HU�~���97���������a���1��2�� L��>�T��<� uj}L��$P��{�'���J쾗��Y��vW���$8� J$��!��$+4vL�5#�Op�a;���c1r��Dqf�ECS$@� t���+z����}_r������.��,. ��ETWג�ｬw�s�=�ܚ1����۫�����2w�� R0>(v�m��W�� ϩ,0WG�VJY�@���vE�K�D����e)*��l+��5��s~Ѫ~d�eOU�C���#�+��(Pp��|��� ��(���� �Bg i�R��ΈD"!3��_y�)�*��� kkk/hK�!UV�ǩOō�Vɢ2���e:?a��'>�Iy�s��F��2XȒ��0�����#�|��z��7����Ϊ��w�:Y=O��j8���m�6�(+���'��0�=ax�6�cQ�{���T�
��Q����nNz*E)g3R��Z�kx�N(�p���h���e���52�W浛�?�U�lT��R\]��v�����&:=�(�\ eKiIJeǵ���n � �0�# �0y6o�$i{}��4�T~!�}��	��ܨ���E�}�,��a�Ltʡ��ҙ�I�\�ZnS
�M�JCʊ�5}��ב`**�V�I�������U��(T��B�%+�8����Ǒ�%�U�BU���!8�`f���O��� ��XhS
cb����>����ʪ�C�����^	�c/_�,��ߐ��q����=2a�2@'��%����̬$"1	�f �r0u3_dq	�I[�����4	�	�L�g�e��[R]�
HU�C>;�	�a�|Vv7�0kY��.�(�����Q���l�Sw��*7"N�	���~<ܔhCبR���F���Efl:���	�ծ1��|�a$�-�׆�n�뫜�����VA����W{}�9����5��;��9�(n�dG\&��2ٟ�T\o���-Ɏ��V�!�PL<��8�6��$���֣�*N�Q �Y���H�� 3EX_G���P�D���>�LS�o5/��ل���`�A:��L.�ZT�����>��7  l�/�5�BA3��*PXƧ��]�r�m�i���ye(�������%���Q��Н��SSS
ēҫ�<;7'��+��KOu���F O$;���iI��m�I!�+�̞�vvs��S5@��5�b>�L�?����d�5�i&������n٧نqݯ�{�S��W(�#,�XD.�a���ֺ�˂2���������S4P	�����cg�-j�~9�e�/b=쵷�y3*��u�^�5���%fWdgcN��-�@O;��9v!O@l�O B�NȦ*���H�d���X�{i�I�NƩa^<�ܑs���b���zOh�k����(�ez)���d��b0!{uA��L�M#䇣�jllTFGF�֍w8�	z��SG�_��;^��<%R�QRV�R -#��s�ŒfV�>
 x������k���ЄBΘ����	
��#
�@��L0j����;z�%��d͋�w�w���kF��� �Tp���K�? e��d~ֻ��~�1|�]7|\0|����ls4l\���軻R4/�t_�F H�,��@�;r�f��+�����\��c�����H�_T��5�y6��׋N��$2���vJo̖��s��4+ɰt��( *��R-֘��BK��Q��Aq� ,�|�v��V����r��=e�z��,���p:� ���X��+H�ܣi|�nU����4 ��g��߯�����T)��Ԑ�0�J���8����kH��'�	2?��@ommU^{�-
GUe��ZE2r���~��i���$�lHY��x�Hb�-e	SQ�zfvVq\I��{
�p�����BQIb��n/�շ�z�ۣ����z���ny � B�%6�z�׽��O�ilk��m����tS�c^�9��٣�c(h��f�O��27�@����y����!���'?+�C��./,��#.ï�k�K{��/lY�ս���؄?�����
�͋74T��6ؐ�xH&�cҧ��ۘ��wY��L+�P<� ��Ug�:+����$<R1��TҐz}mS�M/K���AXO�*�X�Ԟb-�ܦy�h�@��}4 4`����m|@��2;���dt��DB�t�a��N$���ז(�vz)"���`�'���� ��*�oݔX".���N�����g��ܓ
�UN
]���.	*���JH8���)^��+�?~�l)}r�y�(�p�jn�N{��mL�o�Ư�ɓ�9����d�'N<�`6LFޜO1>*�n#�!��
�y ��.//3�����������6A���=G:::�S��,͏J�S��d�=\��:L�����``^�����������^����Ǉ��� RX@��k_��ÜX�T�@4�\_��x����3SP����<�L>C������h�l!�7�� V/��I�dʲ��&��I��b��4NΗ

La�[6����V�z�M��N��8���_����а�c��8��רI6��Ã��,Sh��ޑ����o��1	���җ�o��|
�Q=w6�b��A_�����
���y�����C!�hp������j4)޼,�
���	I�btNb�B���`�J$�S�����o����1]�i���ݕR���Q�Y�>�9/�x�P��9�ŝH��]��p�񩧞b�m}}�r�t&��K��|��}�:yJ&L�bI�x�	��kR���ݸ��X�ʼ�d�P"4giY�f���h�&N�o�}^�LK2� �)#S�ʶ�V���~��9z��<���i���p,�,�Ǯ#�Q�EE�Z�8��!e/�DU��VFI6��8�c�A%h�qJ������Z5���JCBhc�fQ�:33+g������+C��a�|�qyM�<�<c����[oi�E�z��|�����SC�l:-��+2:2J��4T��m�+5:G��yWW�)�*�����s[��CH}&Fx0�� �.@Mqẹp��E���@���)��cz��˂�;�ۦ�cE�޳��l͉�`���<n������?��a����fΦ��++�����2��$�?!���3ʸ;Lu_���o_���]���b��_(�^��A.Gz�Ϣ|o�V�A\p#��DC!�д��}z#�,�e����̍�X�TрZDtj��P,HA��
k�� ����䧬`��I��k��?Hk�׌3���`�׆�[��ա�G	^�����d�G���)�F���~>�^^��կ}]��}��@0��t�y-�LQ��ihp�f&�]226�Ǯ@���b��,��,wY�-�ģ���=�`�^w ��Ĥ�����4�N��S׍�r��
�G�������NV*�5����=~���怅�`Ca�
�8e �^3��6���<������f<I#����dcs�x�ϟg�TA�q��h9�¿ 6{����$_�*�V9��J��K�ع�>�e�j��7y?5�.#��}˯L�.Kz3��U������]6�!�p4�"�Y�Ls�h�!�A����T�Yt$�Xb݃� ����F���PH���/�4��Om � �@0�P@
iR��Ç�#Q�)f2%5�C��ڑ��	��;�ie�%�
���w��19q�;����n(X2š�,����|�@��ٻw�T����0w�R5�(�����$`�S@�u�2�~�4��X�\�c�&��xh룺� -�����7�b��SOȈ>9�Ç���#T$�#!�� �A�<=g��O����u����Ȋ2�o]��_;�"����F�|<�����f[���$�:�E�J�ڏ��[7Y����w�T�ST�U������,۝�Vs�"[?��j͵��pc�.�Y-17BDL�\�0���@KD��S��� ���z��щ0'�4�̱�V��w��r��Gq���se"�a��f��]�n�;C���M�Ѝ��)��#��#�ّ�D*�l����͑��q,`^�
  ��G�ʯ�y �VH��i�G)�:����qT��Ҳܺ�s���_���X�ZXv��ܞ���!�ހܾ}[fg���'��Ç'��ff�dme�����Zm�l���zQ�161��W�&��<v�=z�l6�)����N�@����g@ʉfŜާ�(eǭ�����i�v���ٳg	�n�e:I�6�GWg'Y뷾�t�yY�s�������ia�Y܉c��$����r�6m�Gg9T�6Q�I}��+�ܟ<�#>�3uS3����C����e�/����X7"xo�F����bۡ1VK��n?6 ��"dR
���i����i�!�����q�.F��9eFue@qG5��ַ���Ç���,�>s�n+�b�ȁ4Kroz�X��{T?#�E�'@�Hǎ�wͶ��dldT��mNM����:;.\�,S��L=*��%���+�dyyU:;��	a����T��4��}W��Vep�_��֩��(̱�ue���S�}ү?����w��;��G�����[��F�d�x��#�ÖN����Qӣ �"�>����z�޺=��	6��+�� SD~�{��F0#�PP��J�66��W6�Y׿�y������<�����-v6�+�r|�N�b9 ��'O�\�?i$��#4�x1�ȋbO�E��gw��t��m1Ù!aR�����'��{����'�P�\�ai�.��KD�y�j�j_Ĉ��m�a�u�[���;+`�JuX�����\�zK��_��C��4 6 ��2Q�mBҳ��v��PQ�A)��+�?�峜�:q��R�����m��:L't�տ�d~iURo\���ݕ�u ���\��YW�� �q�\�pI�V7���ix��k=&@����j�������1e�Q�ַr��|�@�4�6��z8�`=�i �#�"�P�f���T�FW�jN_��b��b�	�&���R�����vv��}r��9y�{�k�?-齜��N�!E���nm�Gh�������Z- EX�Vv�s}sG�ʺ;�%�����o�JO�狕C=�2W�A,��ab��VgenyS�V�5���({��S�:�����ݕr�K��3Z�@M��/"�8�M`Q R���2�O�WeYY����P؂0>�JR7��t�B�0W�V��S��_&���4^�� �G0����s/�,���ϲ�t������5�斤~瞼���;�ϳ����1(���q⼗�V�G>y�LOߓ�sr���w(:6�^OH2�*g.�ʖz��Bk?�}:XY�.����p��_w��xN�h{l72 HפX-���kT�G�����#3�>��u���{�k(�_i��Wz���{@A�WYj@L0ŤT�6cfڔ�����qA� ��s��3�����\+ɲ2�����wI��_�����֮t�H��#x��"s��r�츑�o�<��wc��Cq��n)He��at��h2�⊍pZGej`��~�hP�H��|}X���O�P���?�R(�Z@:@�*4�l?�B���e����(�ܔ-�Ñ���$���*"�h@�
d����� �-��9�M�2ւ����� �	yW�u�h���;�H��Ј�x�1P�P�����`�<�я����E�kpp�r��c74:p��<!:t��7���/�� &pL7}NL20��
�~1���Q�;��ek��P���yx��51䪷5� h�}!F%��z�a��iw���#����v�����J- En�a:���������$��#KɆ��Uء�^8u�@���� 6���]����0�7�l��ao�F>�a�Q��4�4(���/a������tȯ�.
H�r�\9��: ��aT����0ˌ~�!e�]�+�H�_����w��K0�)���ˋ��-#ʨ�dvq]�^}GοqI&�������`���ȿ��"ǎ�r�H�}��82g�����s��\e�;;S��)l+�1V�C�?�@�1���cg���h�z�2��0�E�L8Z�疁�#�߷��1ߝ��y�n������3z�t�C`����P(1�U0���h���6#m�GaY�}$����-�0T������T����"��wv����r��my��m�U��D�|��e�H��QL��V湛)K��8�Me�[�����)�K�C�Ro���f�ë��o��{3z=f� �G�8������v�
:8���J5�	��!�4�GMY��T���Ԗ��p�K�4.Q}������d{vwG�pDz��28:)~�i���.�����K�Ց�ѱ.s�#�=�`�!�w��Z���ȃ��n��4�HE�f�y�-MW'�E+�;T07j��[\�5l��+ �U�;����}�C5W%aQ� �i��1UNǘ}����F�}m�ZA�
��x<=Q-wؘ�W{=
�r���D]�i�5S�y�#E�'��ȏB<���������i?!�c��7ޅ�_���o��ڢL�MJG4�Ϣa���8�+K�7��14��ؕK�����~l��r��-�]V�%��⼩�>Ӎ��?�9�Tx�����.F*���ߒ��.y��{k
���7\*����
�Ss���蔂~š[7o��-�ej���/��Q���<�S=#212(O�>��"3woIV�����r��Uy��WehtH��2�{%3ƣ�Qp��V��dl��o4�Ԫ�������_#P��@Ȝ+tp0������C��VaΡ����0�t܁��w��E
�(�M��dS�"������[�p��u�z��3 ���Cu � �i�j�h{=�r嘿X �[����!�����s�_V��(8�d`tB>�7�;�/���l�mI"�Dg���}�zj�E$���`aY�޸'�@L�V���n �S�Te��}6r�^c>�N�(br @@����FS�����[��唑Vi��H���&�ݢ�� d=L�Y�t��I�b2|�#b{�4�F���/F1>d]�FM
��m���o\��o��raOL���ʲ����%�H�nR��h@����m@�?H�6�*C����nܸ+�_M�{'��+�ϹΊ:̱�FΜ��1�02Kv�٦Ì�h�Yl�>�Ɇ�[#�oXn��I 1fĆ?+�>=�|j�ݪ�^��^�γ�p��sA[,������zT��
�9�#xߧ�R�0bnGL�GCb+��G��ܼ�v3r|jR&����S��~�Q�-��1?���7m&��嵴,������}bR��ÀP
��j�*{;����-Wk���;j�G�&u[��)cn҉S'�����<yH�߯��),�>sokfR�|�kv��������y�´�mlK��K�u��v�$L�R,T��෶�%�lZ�^�&[����w���'�2ԅ�T��5�^���Rł�2�B�Y����P*�w4��K&�t�/��˥<�u�.3
�����e8Tv���I�Ӽ��)�Vj�r��9��\*z���}����Z�Isl}�0�U�2�-�r��W�#�a�V�}����^�Z�?���SK�p�=^փRvUo��)Zx��&8�izaKV7�4��a8*=�'��-H	F J�76�4��T��V�+�L�R���A���/)�	h�Zaȣ�tT�L�iȄr,��4y��؛�� ��3HU �Y?��g��~��銴FJת�Y���s�Oh������{�r���%ĲVW0�)@�'���'}�;�n�po��J"����?8(��.�=�}���;�,�G�ޖyR�����ٿ�?�Z����"kˋT`~V��i�`�ܨU�� I48��8��U��XQp:������Tѕ�?.��p�݆
J���{osT]�V�)�8>:{�
ȃ���4+1�S5"��ea{����%VЙ��lG���Ͼ� ��>6��a^A|!/��X��: ���;��l�^�[�k�2�H@����R#���^*���ՐVCe'�z�nM�C�YCĀ�ӕ�uecEI%S�E�I��	�w�I��n+�ԯ�SS$�+�SK�SP�����e��E�A9�ٵe3�f��U3i�VK�^^`{��T�F�QҰ^�dU�c.��//ܓAӉ�!y0?��B�y���}���nV�x�r���Ш����G)�)t�R�sgN���7k��gQ.�.�p �I}��K��Y��IV�!�L���}��Q)xع���)���j��NƢ�ŵ�c����ʆ^��WY̯�3�ѡ����(��-�[��W{}��m^A

rÝ�M����Ѭ���GQ��"b&r4'LZ����@W�&T��L	]ߑ:$2c�M��w��QUk�0JtH�U!��1���y���D�0���ֻ%
,Π���5 |i��@�m��;����ʕ�r��;<#H��K�b�H�x��qm����d;�H$�)~�)� �1*С���*�ܫ
�1��~��Z]Y�* ���w���S2}��lmoI(l�\�X\��v(_*+�u�&/h�.��W�'�$�ҝ�#��6Vuc3��R/�߇ok_7ǫ ?���-�@���������&- 5�<����z��0�[ �ƷL�KƇP��i��IWW�i{�=9~��������-|i��6��ף�,W�Ci ����`�����7���6_��[o��#�Tr��`R���)J*;���^+A��\�J����
�m�WP���[Bt���|�x r�ZuH���,!��z���f�&A)��J����O&���D��/�͗���.+zs�	��(rnB�vP�͛�E�����xCC}�w)3�r��U�K����;�OA;�Q*�1�e��c�859}∌�.�套�'?���<�H4B�dt6A��>�y�bSc��ܹ3�_��� BK�]Y^]ak�#���(Z[+L�?zX��0�6^��z�!��
g@I��pZ�Q��1%q!����i2��^�Sʺ�%�q����7�|����}��2�ǋk�TޟL&COԹ�9�Nble�-j�Gl�,�D5�v�?��.Fj�S�vY! ���:FY�ؽT�0���L��~�+@.#i����P]��~ˢ��"~�Ӛ$�]nU��hl���H������
5�-e�W._�'�8G�|������5�M�'&&��@A�&+�������L����yD�+�,��a}�#��G���П^/g��SO�S
��^>�G� 5$Z�
�����]�{��T��C��۷�)c����\Fh�3�DN�y�Z_�S�O�~�Y���՟d��]y�ߗ����w����#L���q�]0.0Z�L�aƉ�=�7�-���Q���J!��-�ݻw�ǖ��b�7���+o_���u��?�}9s��x�	6;ܕ˘�m1_`��Ќd�}�o���y,�5:k �f5*�������I�i-�Q*����~�>+�`�z��=~��:^u�7}7��lȎf�=]�\Y�yn֠\�lɪ�x�[?H9I�ɹ BR������U9q����ʡ�yj�����&sƨ 
V/}�Ey��y���1<����,L�x��5���%��|����k�nYy�{ddd�Uz0���Cү�
F�_����[.\�"�����\�qCV| �`�pNJ�5|W�;<�-z�<���L��#�B�z���_�����u�"7�\���j�P�)�>��LԴ�68��O��O���b��Gkʀ����uK*�E�g4�x�����_���9�k��9�\ �H���E����_4��L�=�~l��gX�k/�[�r\�ci�q�^\�7E�B��2�_,78��<��Y����`(̫J�52�2:��e^���}V��?+��������d<��z�X9�f���׮]���~[�N�e�``�q����q��*@1G�ѳ���<��'Ȓ=�<+LC`�����겄C~�t���L��|#��h��<!z��^�.����<|�0C�|�`����8q�i	{��@ζY��{��kP��^�� �Ǥsl��'�жi��#EJ�P�ԑ#��*?��lWl�ͧ[��g�kݬ0g���،��>?���(L�:8����w��5�J���מ�e[-�SH��QX�@�5��W�LIA��|��w1R����v`�($��V�J],eg�x��^v���F�S���,dy�$K�xu�57,R
a+��fu�y�͈Á!3�T�*~s�Zs�;._�~M��A��3#'k8T�=�u�L!1-��>��/}�7�	e�О¡l�KC 8H�`*�������W�Wr��U)
�T#��� ����h��n�ٙY����yx�z�f���*�FE�ctccC.^zK�	I�`����H�b���iN�S�Z d� �X��������榾G����b2���n8�X��#���o��7��7/��#M&┐,//�
z��n,!^K����<����^���.����e�[ W3J^8r�}R����NSXm�Z��p�[��6�����6�fz(:b��0fN�A�=����6Y��}��!{M?��HM$ ƳE4dZ!UX @��XЂ���dO� ���'O���3�Kg�s��}UCYT�C4H���8=-�F]�tI.�yAL�_�s�+� ?��֋bL�bf>�� ��2}���ȫ���I�f���+�ב�	X]
>a����i0R�Ѝ�2x�6�m�x����_��vV�z�In/���dһ�}XV���-�*
�Q�È(k��Fۆq�]��4̠�U=��{��=�����a��
-/�z ����OC^?��<�����c2>6BS�����K�������@��ƌ���:V���ף��8��P8a�y���b�����t�8�)`\g�i@�A mv�[�#`��Bo�x܌U�Mm�&�}�J�6M�3*� &��Ӵ�r������ �B&��C��)o�Rc����ٟ����R�ds��)�j��@^���q��=C�nz{w[�߸./��}Y[[�/|�K�4�@p=t��0Ä�S�^0^ӭ�R��t�g�А|��ͥ�����i����ۿ�Ϲ�qR.���b��6����ǟ�x"���\���G9����I�P��Νy�v�9c6UݸB�(��(���B*�o��1�0�[��V�,�
��fCy����a�z#����f�A�'��299!ʖ�~��r��hy��F���X������B�T���G���7z䡍X%��\3�0#�29ӖYF�@m�k�/���#���;���#)Z�hDE�;o�g��#Bo�7�C��6tI�eQ��b!��������A3U3�~� pFF��w�KGg�䕙��VV���U�i��esywZ�G�NM�.����C��i�291A��ZՑKo]R&�'[[�t���n���sVj���G����༩�tIf��9޺�����-����k"��n�
ݷ�l�3DΘ4�5v�0C}|����$P"������:� Q|cH��Ǵ��fZ%��vz�#a�|��9�ev�Ģ!2k��>�6%m�Gf��.�5�+-W���'~n��m��W���0g[�c����j�e��R������>�����wQ�q�5Y��ܠ�`ʸ �m7C�<���n��Ջz�������̕��#�[M�����G�"cѸ��{�,��e6��/��������c�R&��㫺��hX<d�ZŸ����?/�N����5�y�&�� H�,Wf�=��ϋQ#�ݼ"Ejv�I�1��Va�lH(�aX1�e�d��?��eF1���<�1�<*������Q/Ƈ6|�	X~��N�� ��H��U�~��9�Y�:0����Ɩ�����@%qP3����n�H��QX@&v�9ӓ��m0����y�V�=�:+.4)���.nʽ)����Ҟ"/�5��~(��ݻ��z��Q6�u6�E��p�'C��R0�mYY��dQ����l�y�檻�2��#LG�@�޽���g�ַ�#�<�Aj`hH��"��0�s�3��y�1e�~t��"��������]=�ޗ�^;O��3vF�u�G�Z8W�M��ED�$EL.hJ0P6��������L�_����FǓ��u�t�������/ ���>׺�g>o������%��1j�9��N�)R}�+���.}?Jl���6�-!m�Gl5���;H�v�dt��?�2@���ij5��n5g̓�6�K56���[�"�ڔ�62>�_�S7_�p2��K?�H�	Uٗ&x��z�7��{x}��ȑm�W^���(K0���䉓r��ie~��u��C
TmWw���
s����������_���1�엁�~vElnn�c�21>!=�=
�hʟ>y����9e���]��!}�T�X,Io��w�yIL�0�nH���8Gm��0��hk���Z,������Å)
��u��l~����(-�`yg! �DzT0u=a7���f�T�x�0E!O��T�Ƽ��Q0�����.W;�{kp��� �2�?�d��Zn'�e��Ey�cjT�ф��3gj$7��h)�j�Ж�Im�I3�w;�̷��R[	��$����nB�Q����#�~��r����ɇ>�q9v�����%��/2��  E2�b5� lȹBT{��]9}�E�����n�/���?D�׮_��׮�m�Ϟ9#�6�k�`fV�GK4��l6#++Y��Fj��X�Q�n�< �ܾmZg=ޖ8�#�4�����	�>p�·y4�y�8`h��S����ml0��v���^*���8��X3�S���Q0>���+�6	�3�x,��p(r������G)Mjڴ���E	��UD�;�;L��{�Ӄ(V�؄�� -��YIOO�l����4C)���7"O�A0�"��V��f�Z�%[ȿO��:�`����I�v���`�� �<w�	9�`������������D�������?��:U.+�B������|����M"d�Lx�w�lE�#
�gN�d����GV�g/��lt���f��z�<8*###�DHQ)o�s�9�x���`y5�#Z*�����A��NN�Tx� NH�8����L(C���c���-H�PH�sֽe,��	�¢��ȷ2\��5�V��l��y�����o��Omm�Gg5��X�Go��Цje{{[��/������B0��˛׃&h�D�k��) �UR�S`�9��H��V�ޭW��ߢ�M�w�"d�־�ѕ@����c��F9_�NT�Ɏ��6�u��1�:x��5���d�6�����7$]]�l+]^Y����L�����](䔱�HWgJ�b�SW���S L(�CY]�_�'�`T�z��ޠ�5~�i�bN�[8h@�lq^ݮp\�*�4F�U���&�DN`_P�Qq��7/�87BSD���B-V���*��bP��P�I3 ����ٺ�B7I���QztwuHG*A� �d��Fh�ګ��e��48����5�'�3�����7{���Q�E�q�U�����d������Ӡ���u�ɡ�w�ϏP��K�>��I	��,',���`P���G���7�l�
���s%w4G��� ��PC3���칧d��]�{oN�:���q�t��D���3$[���{	R�;����htpD/����2����3�N�&�׃��C�֟e�嗾'����ԓ�Ç�˃�E�/����u�>W�VO@z��eecC�7�2������~�dltL��$���Wߔ�<�]	)KE�B�F/�\�Q� Xw*��$�J��BQ8� �``l��Rb�),��
v�|�je�>����	�i��(ZG��#��*R)�|���W��⽌m��f�0��(�/��]���*��Rn]����	�J����]hbm̶��j�Gc� �fT;	^�L�u�B:�څ�y���G>\�8P%#���uP�-S�͠:���`��~Ԫ%:�7�j)�*E�@aꋜY��� �z�����Bb��S�̌8A���#���wZ��M�!jS��*���~}���R��C�O<#���w�/��+�.�c=���O�k	��H`GJ���[	��u|��Wd7����M髧����1(��.����'�̙'eiqC�߼/�����ɹ'?$�i���H�Tٙ/'������˖���!��\�v[A{Y���ܸ~]�O@&Lʵ�WhB�0t]��3�҇���Y�t�2߉�T�j�3��Ae�A���8���st2��|ܴʒ���k��T<���h<�|v[��<�� ����1Ix=�Ź����ewWx�G/�5/�^�2:�-�C�����uߕM�(ә�j�_�rZ�!S�n�����p�P]�^��g�ԑVQ�E�P��9�v(������06�}\%���m�p@"���,�C�,����)�2zc5$K�&�!5�8ڂ�j�8
 (Zl7?�V.��V6���
p����t�*��\���������_��rv��j��Ѧ�.F5ӱ�x5��Ǖ�&��Hv�H���lo���ޮ|�P�'?|R�7��|$��_$� <6%�·���[2;��!BA^z�U�����f5�ϭ�M���ޓ+����A"t��!	�5��=�|#S ����E7(� C!Ț�Ek�o9A^���3'�$J�br�NDߛ��m���v��k��-;vLfK������tyB=���49�O���m���C�ҍ)��j
���X�}��j�v�F��)r�S��!��}�<)���e���>?e6k3/f5����Pd�z�`�%�]}��G��Dq	y��A���*�S������M���(d{mI�
X>r����cK��#��(M����JLъ�E��[��G� ����xL>����mrff��w�v0/� ��>�%e�1e�	}��f4\v�b���/W%]h�G�k"�c��������5�r��t��������o���Ш�4��,Ԉ����V�����da~���CC�1B٥tSY^N�iKY�6u��XT:S́�
 �̤��_���!��ݝnл��q:L����'.�ݓ�.�ۿ�W,O>�$Y�ݻw��6Xt�!\(��}�1���.�����e�'b�zq}n/M�gg�8��m4{m0m�Ga5�>=��4�N��_1d~f m��2_DgeA^Aj�QvRٓ�U_OT���drl�y3�]��vV�TKR����7�D�+eR�������d�H��?�ASf�xx�<1���_���յ�á�P$n��6�����Ɛ�E�szJ���H
4}�1	�!ܠ�9�JE�\S��W������_�������L=ܸ�(�r26%I���\�:/����p�<v����e�j*���/9���5uT̑���}�����0I+�H���g?����gqI7�P !�h����	�ۺ!䙣�Wd�(�����@�$��l���ط2�0ˈ
���̯<#O�{B���dc}C�;(�z��ӝ����q6ԁɃ̓����3���ܐ>���ƺt����63������Q]����g�NQ�]^Z���z~�EF
��90�|P݅1��@�E��G�ɉ�1�M����6'��s�����>D�^�񊲩�甆��I�L�df~E������A���2�g���2l�b *>l�����κG<1�E��OJ8f��ɐ9~�@�:�⩘���I�YGX����&7w�����ޡ!��[��~E���EB&UPp���eY[Z���q}�Y]_Q���S'O����(�T��M��* !�H��!Ǝ���e�c�9뛽G"�	=<)5�O$u#Pf8�0'��<:�ّ��wwW�tu�p���nF2{�zm*ʲm��Hw,�_��Yd��g~M:�\F�{��w�W^��|��r��9�T�y��\���ɟ�7��ɂ�׷��;7t{�c^__���AZ��㡚@jۦj�&���(�f��!-W�n��Qv͌w��EH�ʽR�()��*�V�"�RY"~K�G���TP��m��ٻ��x_Cд���D�[��8���[���!���fX��R�H:_��-KUCI ���9�הe)�������?���(�tw�iH�Ņy��?#�� ��c�-2@[^!2�=&@��]�`� SG���+:��	�1�wv����LϮ��wf�����$�'�>"��=��pBd�`�h۵��JY��1�y(S��6�G����'�Ͽ&��=r���$�Q�+��-�C����������an�|�xֶ�܀B�|a0¶O}c;tC{��1��Ʉ�&1�X[Y��Ug%��EB�;�f/\x���Y�&��A9$T:描��{B����Ӫ������Xtb[t����M����O�������S�4��h�6�<*��<��9>5!���V�f��ͫ����a~BN�>%�=�5dE��0�0(�+r���l)���f�II}yGʸ�KE�4[LW�|EM�����)*�5N-Hwg��+�u����%�MH�R�8���h
��ˠ��.��lР�u��L&'�o������I��W|%�}��,�!�K E4�x&��p�[��
�0"y������+p�еV�="GJ�~�tUW��<#R_���$�����elr\^;^�ߺ&E��9~�	�|w�GG)�����W9����$
Y��h����?G�Ba���x��ɓ�	���y\¡m �0�5ԇp��ۡ��f_�~�a�1��ʻ��ګ�>�e�1�ƾu�ސ3F	)8�JA0���~fJ ��'���^��c�PWRN԰�W2��2��mɥ�v�CS�������� ���!'&p�`^���!�ܝ����U��l�6�RŊۻ��l
h0�H�CR�奠��Qd7�m4�_[Oԧ��%�l������2�tF���}]ң��&�3pC��.d����&����:{��Bg�s�s�o!�˧�R-��g�c�%�'/V�z��+@��CT�/���|�k_���>C �RV�B�>��!��m�#N��a[�)�	=����K/��ῐ�|�3�������i3��;*�N�uY��@����=�xN�F�M�%�z�=����|oݚ�c����G��i���{/�.w�ܕ��#������_�/��V�>7�衳���3j˵k7�cF��ɓ��_��4�ٵW{�<��}ݔ�Â���� �q�=���@���){���ba1j	�w�G��Ů�e��ݑ������z���-*UT����:���ܤ�7�_�cR�ȀlomJ$��R���f���:��R^Q����v9��1��hi%�HR���ٕ[�o��Ύ|�#O���'ex�S�!,U(�5m�Ln�8�C��ɡ&�l��=v@�A���_�7.�I�+�?W0�lHOU��n��
%e�6��1�ޡT���26:,����-�c���Ds�P��H_�0��0�v��^[$D����JgW�ܹ�z٣Ǐˡ#��I����[8UEeiyM�kL����7���yZDwYx���������.I,~Wvw���3r���>�N��ƌIIH<3����E�����Δ<��9�����>����h��c��^����f�z�ڏ�����,��qfBM���?��Z-��J�@�5��}2��)	e8�sӒS�t��)9�x���Eeu
��W�a�#!۸��C�Y��;{Fo«����as\_�"Ё�Vk�ݽP(�k��<��z�i2�p����;�B������1M��C(��_S�W����l��C�o�m����i�(zk�,��+�4wOaX��Q�"A��ʎ벛�U���檪l2�k�W���~[�Fz�i��߼yC�u3��7_�p3�KRݤL'��`��2�H�S�!%+(;{e�.n���,��1�٩;'����0�ϑ1�y�>�<���� ̸Z��ҕw謏���ʉ7�U}.8U����+(��_��L_-�)�BWܦ wBQ������Ye�O>�D���l-���^I��c�e{�J��݀t��i�Mx	
`Z��!�����t$br���$,&a@Z,V@	��4*�����yN�L���'���U6��5\�h��T�.D͛�i{G1�b��07��71Xon���s��ܞ��MI��
�1�u�|����Cu�δ�N�Q��8�8k��4���zN�b��֊�Ir\�|��������2>>���T r�>/� �L5�H�e_���4�u��LNN�w����y���F��������f,�l.����ˠ��7?C@F�ԝF3��HC������tx�{�`-�t3���ާ��!��,1�U�/,ɔW�D�M�x���{�{EnpL��*dø��A~��^���?kK�W��@���d�R)�B���>ʏ�>K1�ﱤ�ۓ���.{���2���u$ �9@�����:N��������q��ON�>%o�}[֕	�J{KU�m_��Jd36��0��Α��9��5��L6C���C�����K������".\ԝ%���g>}�0/p#<5.0�hçSY���p|���X<�K�"h �dF�#ю�4t)���G�R^�pX&Fe��=�ދ��巯0}������#,��'�?�hiRh�>��g�ԩӒ�HJV��׿�mIu���踤�f�y6;,//ф��uJI��^2�0�@�b�$^}C`X���ð��vކ��R������S_�I�^� �t���W���{�2(�I��R�����1��D�	2�z����l ��	��^��2���!�� B���cs�O����=v�[4��6�!�G��\`&�Ǽ^8D�ʂ�zwz�T�o��!�'���=���0G��/HWLe"NT����}
v�ˎ%����f����!h0ԟWx��$+z<{۫RP���ө�c^�00?����6�qU���{̘��-�t����2�<b>�X�(��)�����NM7�D BQ}![� ?��|a�Ϧi�����*��)��'�&�)YX\��a�!���z�ȡ�G�_��?�,4#��W|�N���x7B��J^�8���7��m�'ݗ�߳M���r�I��9B6? d�b�
�<�=��0��/�m\��2GA7�0L����s,�+,K<1-��^�mQ~{�r-��L��)��677�8�3j�ǮV��U�`����>����ڲL߿�?���K@ӄ�N�<���Ao��ȀO��]8u�xnno*���hP�6��üf �����p@*�m�y�a��������\Vbɸ2�A1����7�O?{FΜz��08���R,�,.����G��L:�����^��_{C�xC�ɦ��mwg�`
�fM/��vZ�7v���X�A����G����C�`�P<t�0���Ҋ�P���O>F���/�����Sf�����]���$H#�j���������� �@0���c�=�� Q�qha��וi�� �5F�@����UL�P�qL��C��i��!���M+.6=/��	\�Bhx��	N�x������5*
t�}{�2-��o�j��˲xo��L���];����&dtL�!hggR�o*@�I
Bxe(��c�Ž11K"s�.h��	����͛=�$�dGS0�U^NN���4�JJ>�=�}SY���R+�0a�_����TW�`
 )KM%z%�JOW����+k*j(^�s�M���G�LM)�*��ܜ�����\|����HY�*�ڑ��t��W+�����+�!�� 7���ʜ�����s�W�+�ܖ��'Ȃ12�b�Lv�V���1�����^?O�/���X 2>�zΥ�C������P�10�C���Z ?���'E~j!�.1�1��� Mѱc�,����~��F��3����\ ��]��(���)ړq���Fa�m0m�_��5�x�:�ʏ����O�ԑ*��� ��/9��W��>1#=
��ؽ���+�����Tq ��̍F����y�@@¡�d�5Y����K�ބ齬�
0
��B�H��ƭ�
R�d$�'�^���Cc�����e949%
��Ǚ�q�Eq5�HWw��ݹ+�3�hg���"�]][��׮J*�@P\X�հ�/���O�#���2�����[�nq��G���2�AYY^�������/O7�]YZ^�[�o��Ɔ<v�d����K%�����Cz>]2;;/�̮�(zh|(䲬�WؠP# B&5�E�z}n��>�h�R��#�b;U�|����;���b���Z���a ��a���D�E�nj����f�="	����;u@�O��P$��n��ޔ�%�=�KH�z�g{�����~����!�ć�g�2�9�M������pB��c������3�=L��M�bՒ��LEbCz�4dyeIGF$
;�(u��~�><u�J���Y@�q���y�m��eWkpjH(�H	yGŎ����ݴ���H�#3��1V��Xĕ1�o{G�,�Ǟ8A �k�mn��щ �~zX4�p+�Y��0J ����J� �]1���|L&'�鐟J%������㣃��s��e�ʁ�a9~tJ�|�ڋ��U�C��؈�o�+�d���k�H�\��
�I���e�\_V�<L E��7&$ Q���c���zS���?��(+��]++�:'У�\![Ŏj���,���RZ���=�K�E�' �a�l�q���	i$�ίzͤ:h�U���~��{w�P*(���~��A*�m��^���� ����f�o�@A�Œ�n=��> �?`4�jQ��*6�4^\Y�ա$g$�:�egcQ��6dp(@�����(2P��n��!�\ߖ7�_�+��v��n�m���ĥr�]�+�A��<v	����O�������s�����V���=�P`Xb���v������3�ȏ=����1�	�Ywvw�H������P���5�@q*�P��!���ܹs_�?.[ƣ`�THOoY����t��u��W_��.]��ϝ���a�YYY�.��������-î	g
�u�1�X�dt��]W
�P�K��9���<y�KȄ�uw�v��ձ�vs蛆�J��~�0��ț�o���K�Sq'�*cU�ꆳ�U�ۍ�������_�����?u�na�d��
���1���˰,3K�x��-��i�%a���P��[���*�Εk�������<6�'���=�}�.M2����u�:�u��a�d $�D����<X���ue`���]��p͑����B�a���l��w�eP�YN�\!�3ZUcuM�?Ʈ�����N�(ǭ�[���`a��,���I� ̮���윬��8��8�����mm��x]�)���p]�{L�����a�ב���1'׮^�ٹy2CtO /i����6�e��4jѣd�p��[U��WKy~��$�1���D��Ӧ�˶�]��.��Dq}��=/r�� '�����U������jE�}sx^��a��\ڑF93����]�yQ�7�i��h���%X�K43 �݇�攐��paaA6��z��TW �Ӻޔ��'{��<X^�~{]����ٙY��/)	�ӒGoD�39̪ވ!�
��rof�,m�������#�L�E�� �F�$4��ժ&�cz����&$!Q�Ҡ�?88��]s���� �?����#���%� {n�Y�ˤ[�2<������N���g	V����.�̻���������255%�?���;����XQv<�����6����0���|�K�=D���$��5۔͵5��a���M��\���sTK�\?�n�5�6�3���1��366&]]]�y����P��g�l����两�)�g��A�?:2�@:.��������-e�n~h�`U�ji{���M@�-�y�y�c�����9�\{6�hH/M���EHC���=�]\�1e㇎i�< �[�͗dA5�CWQ��Tg���9YZ^��Wo��ڶ��q�b��xK*��~�5BJ����H�p�CDn*��gf�h�=��n&��0�Hutr�p\�`�esC٣O�PХ8�]l �x̸�Hl�+�����R.�'��I,cu���d�gN�!�q  ��?�g��ѭ��w~�weJ�|&��9e�����I<���3sd����}����4��Gvo]v���V�IL����C츀X"�
���\#�����;����~�az�:9�����������C&��eJ@�9�`:I���(�=rX�#*+ˋr��Ρ�X!n�mק���\��IsW(c�/������f��[fԈ~�5̵m?u�
k
�5Ҍ\�5� �'g���ã�N�dK��g�ݐ�ަd
ʔE	�|R��^0&�N�YBַ2�l�����v.����S�xHCf� G�
iN�h%�'�%�,L20VĻ�7@p��U=@[:�����h�8����!Ƽ�	@ �Hcs�c2:<$=�
1:P�lo*�\���V��=xz���1�� �
NȽZ�Sgq��֭wFc�3dT �=e�!��0��5����&+K��6��=-�b�~llTN>v���� (����$���0^fZ����6Uo~��f���
���Fu�$+���/}��:���b���rQ�7B#ꊲ���������ӄC5���n�i{��,��䶱��f`])0����MN� �0��^���P\�5B��S܋3���+��=��ڑ����P/�=(qW�GW
���-��X�G����=T�܃U��d�\Y��}�7�*>��0LNY���3%#A�涌�z�n{�yO�X9#��4Z\�;�`�s��M�yCb7 ]L(.�����5������C�;<4�����n�����|ꓟ�=�GNC�:g�lR�ڸ�ʥb��+W.ˠ>VVV����ttv�c���b�}�ew�=Ǯ4�:A~���&g�>#����r��Y�\_����8?-�Ї��r��u���g�s��'�r� ��\�S�Q��6�
з�Ǥw7d~���ԉ#lu]Y���^|^���/J_�a���'7 +@Կ�]fȎ�K�2)��1���*�FN���6�ۅ����Z� q�x�7M�%�뢠��*j�s�����ߎ[�ݯ�3�"���sZ%�.�����
�,;�ľ{�geVU�7m�ݴ�0 �+���+�R�$J��*҃�/
��I�z�BzTl�jEjI�@� 	7� ���������^��ι�fUu��3� �}����ʼ��{����~/=�0%Yu����e�`������Xn�t�b՚��+�h4��δ����eq��}�ʈ�Ny�LN��_^�`jw���.FJy�7�ymI�q
�5������\U�����`�V���������� ����e�>]m�V���fKKwČ����I���,��;whN��q��M���i��u�y<��sX�Z�o�)�X��Ʀ�U����G����(�����g�Ǐ~�c���;*$BmR����d�����������3z���;�w�{c#�8}�^����~�" �(�2A�!��1�&��d�rK� 9�=��Ҙ���rg2�����G"J����濽U���f.��:���b~@�=��[wZ���>���es6��Y�K�W��FwqqaQ��'N��M�_&[����0�����]��	�u�sCJ�j�6P[����ed>��� a�@
���)(Q��hi���J��+E�cz$��é��m�H�*3&�1�mT�J��nT�c*rH��D���.kh��Y�8����[�����̴r-	�����J�}hpX�Y��3�Ca�7_}U�e[[M���UN��s�^����XXXR��))(����o�s���ܒ��'���E�Mc�e�|�7���V(W7��)�V����rZ��ۤ\���W�*��2��z�i]%��[ۛ8) Ka����y��-i�v�`: �<y�r�d`w^���9�:����4�m?�V���a�.�r�K�A�C}�kT�����@z�����ƍ�=	��z�4JXy��M�����vpJӖ�/ϾmbDq䐵Ӧ�	��%�i~9��T3���nS��2�
@ix�^@+�Wn"�9ir8��;�*SZ��������1���D�Q�$49�/��&VmN�VhVW��Z��5����g<�I�+W�aaqǏ�Pn����WZ�⪳C��Q._D�]GU��� ��ڊ��Z�H��1Y�g?�mc�lv�����$2�A���kJ�}L��n����=W��;��7���s���{k�^VU �-���K7��?�.F�اN�R ;�*Ν����,ad|Z�l��eL	��8��1��3�Q&�t11��ƫ��%r-�����?��鴻����Wp�Ƃ���U�	p���xB�٧�zRɬ�o�N/=������S�)6��t�Wu����ggDF��"�&�4q����O��^F����3^i8�a�a(70q9������W�άXq�˞Ho':,�ӳ��I��h,u'yQ�&XHW�T����*(1q���\�|E/�����^�;x��M��H�g�<1
�����#�(��I���b�<� ��	uC� �=��y|����v�%����%)�|��5�;w^;m20�����;
�G�W���u�y��.��W,O��
�d����H���>�6��7e��ү~�f��F�����jK�F�i�6�b<S�&�K,��X�YQ�Jh*ovyuE�t��~���e94{��o
��fc����������P5I}ՊMkrK����~W��ۧi3*���dd���Yr�`5:��R���kQ?�A)�$I7��iy��)��C�~�Y�^Ϸ$������bb̸�>�v�0I�؟��Xs�P=�P��L:���f&��b#�_�������o��_+��>-&��\]�~M�q�F$�����a����N?��}�Q36�͔���+3��O_��~�3�l4�jI%�2)��*7�������j�����9�mq�ocP,e���h{����C�Cn`'��0Ǐ~�*^@�{~P��'���["�2sΌ=+������)��vm[9���7����E�SX�dҙ�a�܇W|����YU����z�=�E�<�U�Ǝx$\h4��dY:kS�#���S�A���8c�acc]��{��|w��<T���i��*˿d��dS���@�{���Oi}8A�pBs�g����l�g��M�	4=���Y 5��v�E=�P����X���3Y�{��{���U|�[��$K1�Z�Ӎ�F��?��!-��{�s��9���(g���MzVMɊĠ88���4��^Ç��`��kx	��UԷV0P�*��=�1,�Ӆ�`JŦ�B����I%���y�4ַ�����+��1�~{���r�MMt���b��=��ݶR9���Ji�)�a��b*j������-����Ҳz��+EY\Z�quh�$��!@\S��@	O<��;*�DMuaS=φ_B�6������Ӱ.�盎�]��eꪾ�c�*����!s�L����׼��x�a�Yt����+�)���)+�kz5��A=��	Mne��g=�MWO�K�Q�i��-6�x�JķY5Zb���u��/}Y�N�%Hj���(�	c�9K��+���k׮��R�2VF;�`y��WY�ɯ������_\Ge� ��P�cq��ѡa��dqhk��8P��PҾX�9**��= o,Uq�f�*v�YZx9l�;(�(��W �u�8�@� WQ�=�T6�c�Z���C+vMk�e�b�u��Im�^F<�-����s�{�i���S��F����k�U7�# �w��u��TR9E_�[� �3t`"�����O�����1i������"UkHCWiSʬ-�.^�6�l"�k[�K=�g{�k�U�ۛ�����<[C�D�i]ۙS�S6��Z���X\5١�����%<�gD���x0��z�is�T��1K&����_�����O����_]�s/�ո�r�$�[������;J��B�����������C�&Ю��t"�$���J^\�@!萡ЕEk[\q�U)�L\]��wT��� ��dC�_����4X*�<4�EL�QM�w!�D��5}���R��&YI�7���j�wjZ�5�)�e��V���@�˷U��r�����\��K_�
�&*x㵗q��U�����Z����{�]@�_"z�4l�-3��>��{z�Ϧ���%���V(�%��*��f��j�!�I)J�v�dW��]��CϾgrH���N�DŅCDqQ�9D�<����LStZ[�0���q���<��޼4��#.s�C�J��mV��~D��A�lD~x��YL��j�o�����X7�ҝ��`���c��i�Wt���8�����E���Xp��k��V�FPm��Sz�R&��	!̋ś-���'�K���ۨ2a�%c���\N�I�4�rDk5�uu9��)���
�&�x�l����V{�PF� ���z�j�k����Y���4C��������b��^�ыx睷taZZZ�c��}Q'���t#�|?Fz��l)�SO9�@�q���fJD}6�3N���֏���T�2���N9|W_^��I�4-Kk��I���jSh�1�I����Q��@7��)PK�{���P�3W�ϖ�I��?~���17SA9+V��1QU�?*�=�LXZτ|T��rT���-���7qua�s�0��7k�}���S��2����*��YU�i��j�R��9,n����ѣ�K��.K+�͓-X�=�r�Kkb��ə�^�x�X���k7�(apbR� UVf���W���2��EI�x��WY�)��������R����t��Ԇ{P(��*OZ����m���E3f�CR��&�d付����O�1�O�z���159�m��i۷�IE��C܏���>%�#�����GX���C	*J69j��东��Җ|�o3�N<Ib?r����U��ㇺ�����j�:�0�2,Mv	�o�X�8t��\������qpF��a�t`�Ff�
8 �uF%�y�kJLogJ�����m�R����X�YqХfM��� eK+���|���q������>�������4�kձt��0�M���Ǿ�p[\�A}��[�`u��o����k�cl��b�u�j5T����!�I@@=�e�4���JeP�j��>S����M�4I�>Pa��n4Z(�e�����xf��e�-�*�i��% ��@�ZД;$�i8�iq��4��3 s����oQ��&��-⑺i���5i�A7{Ьl�@�3�M�:>v�]�3�o������]�jyF�ʷ�ҳQS��8c�*>)1_,��	l�.����ak}Mc���+����D�BF���D�I`d����8�Ņn���J�TU��nj���}V#ն�ڣ�Ϧ��Y.�)����Ϳ�w��G8y� �\��������}'O�Ѿ����/p��r�Q9�o/,��7�A��T�P�`*#c
�#b���p�&�n���cp�����3v�%�Q�^u	z=�gMe�2FY�d�z�ã�30!�@�d�z�j����h�x/k&]����#7��@�JjxG[����o��-��8Jҿ��x�:K��lQD������[�$	��Hϱ�
D�����5=����*6�4����P��L��U�J��"��-$c��n`H��[i�2^K�:]�t>���5��ZD@������@㓬d`�Z�����tj��]�����W����Ν�� ��}
����N�>���<��������^��X�7/	@5Q���eT5�nm�`�8�S�����Ё�:���9{�]��ʛ8r�(�y�1�vזW�Wt!8|�8��aqmo�{�U`�L=��t�x*�Ga�vK�X��i场��N��u��ג�Q*�Ժ��޲���7I����ۧcs�c	����-F��O���o p�焂���	W�s�Ha�uJa��?�P�oEU�ah3���5�G:�'�=�D�@3��erb!���҄4�f���^U��ݖ�d�5�
�(w��m���Q�75
F��������i/%��P��84���� MZ�6f̏�:�3S��7�	�W��<������'�0ԬqÙ�<~�7���$ccSx�70Rǳ�}_����3��Sx�g���op��,^o�K��/<���wO>>�<���+��7�������?Ge���Ml�l2���Y��xx�l�1?V�h��]�4N��S���j�hkm�X���!�1�&����8>$'Ӽ�����+|��}�6�������h{� ��֍:�<�"	��(*�L_��ǎ�D@�T�����ht��狵�t%J��em4kz~-�w�Z�ϵc��0�U	���
!_lHy��律�@ɋ����5�CХeKk�@Ks�z�tW��M�V[����l�Ǉ�/������k����wq`ʴGn5�)FRʀu
�=� ��ƛo�#`Ie�C��1�c�x��q��`?��z�_����������DV�|�3��Ye���m��eL�ajP@���
О�[kZ�Ī$R��͎Z�hw���h�'�L"�?ebԡV����e�g9u���j?֍�.V0�i{/�����/��yD��	JgbK;��o��q���*:�3�>�5���6���dVk5���_v�#���0�=/�aK9�`u��u���A���B�,g�|���R���o�|ri��]o5,���-s@�����^��fw�3�h2�%��vӨ[�g.�������&&���[j87�آ��|����sO����;���w���9�
Y=��J'����8u�(~�׾��sS�k�Z5\�|&�#��p�.��?=9��[v0�: �\�͛u���+ڃ��H��
4�ܻ00U�^c�E��2
̵�-S�877�L�����sF�K,����ۧdK��1��%�� �e�V�٣@j����.��[�왗~?0ɣ�&�,�n⼒�l�7ʌy~�u ύn9���R�LN��U	�ߓ	��;\�)�~D�x���s��x���&t�zb	)+��5�r�@@P[�������𐶭f�ۧ�x���?� �R^(]zv M�����K��Ҳp��W���S|�{���?��8^��fUK3}�9q��*����2�����"�����*�����x�����*Q�(fm���+7o���3|���B��2yH]�f�e�MʆOz���Ӣ��_.�*��=8,�eo*~C�U��X����7E�o��-�U���]��%V�P�*����픧��2�	�T^/��i���tZ����q��� l<�BQ���}�3���h��CW�XH|Y:��J8F^������`?i9��&��ҥ��	�Z�3�ߴ�S`
��)��|9/�nW���Պe,�]3M�HJ�Ccae3i1��<���;�qل.��Q����F~bf�o�ccm�SX�1Q���p��GU܃J�/��:��2��������]��=8��_�9���o�K_xS���BS���r��A�Ĥ���-�ٟ}ǎQ e�<PKKz�>1����W^�9����/��e���=��6�-KY�����)���5�Vi_�P� �^���g��d���K��������3��_��&����T�����ۧf#&���0�Q�0?���Fɦ��m/-M��o5��Ҭ��?O��tE��XB��R�b1+@�S7��?ڴN��@¶LFr!{ͺ
cd��Vw��� �ٳ��'�ۮ�Bs�3gaԟ��c����:�Z��)���Z����t�*S����˧�jh[;sQ��vJ��(T-g���g<�g�A�F#��	��L���w��>�ҝ-LW��g��?���v�L�_����w��00�͵MdC���S��=y��BJ��Y��F{)��]����;)���SN�����BQ(P,`rz� ����zMij)�H�9�=e[���CU��Y*��k���s1�%����*D=T.�{#�I����w���]�HiM�;�hb2vHk��M���BskAs[\b�ne��� �d��IF��K�����X�5Q�`eTA�-�d6/�c�X�������������W���iQ�D,��&�Hi"(���Z4@�L-}�O���3֗�)D	�{�c�-jê$`�v����{YP��-��y�ł�
�z��(a⁇��\�[�j_;�:9u���_�D�ir��\YD� h~c��f�bi~E�C�_2�5�3���� g�:�ɶ̔A �5X�S�X�My�-��GGph�0�fgp���=/���tn@�LaTIq���g+��*u�s��+�S���5[.�>uZ<�:��6՚�gӆ�v�,����H&c|�|JNN8fvӡL*�(����513=��c�055�]3;�.]8�u��4�����a\�rC��h�104���N}[-Ĕ#�%�<F&~�&�ri(�uU��c��0��&9>V�#��_��
��ː*�����^ߦ$]S�=�o��69��-�|�$����
ǧ$��PY^C���lnU�ڧ<} ӳ�QΊ��k�۝} ʩ��r�8GP�����O�X{J�O�0�x�����gy��R���_�N�L�1$�k���srW�=��'O���/�έ[8x�Am��%�u��h��-�PF�h��ÈX��g�{N�ta�nܸbx�>L,�>�����m�lj�,�1;K��]��Q]3h'�fp��$��CehX������%�����<��_C�2���x�X^��El	��(�����Z��k�T���Q�,A�ש��<A�'hX���-���2h4�� �����\�����n��������P.%�w��^A�����dm-K4)α�����Ul-�cu�'@:���#�`�G3����"2���VO��գ����n�S�_�Sk�P�񩩞i!���u��FP,���[�b�p��1��?�9��X�%�on`��m-�,tL�6���|_�����˸x�&�pac���R�e����r��R�/���wߓ�]���k�z��*cgtp�����L�;ZjT�f�׵ɇ�vě`��gpznJ	O��k�q����.:1��O����e\�|��\@el
��x3���XY�j��G��MG_�论�=Y�S J�k� i9�����S
�XY�i���O�]�(0��,akm��6�~���L���d��G:ø`��LlꆐV,I�Y=0���� �r�:���C|������1y`�PB�UE(�����3�z�ŋA��*�����T�\�ԇ��x��04\B��V��S���O?�J���ǎ�0>�/�KjI�JEm�GMֹ#sZm�� lL�7�T}�a���������X����i���B"I��]�ll�(�m�m;2Ve1a�+��bߤ@��6%�Q���wo�j�i���=r)��N���3�qxv��qobsm]��P1��q�:1'.�� �.�����¥�X�}A���2�3� �FI���2��	q��W�V�g�La1��:��%mi�PWAP)K�<3�D��vC�x��E�:ۘ-��䈾�t�u��e,��`C�6Ry�"(�f~ �(.�!<(`721�G�O�СI������,W/h{�C'Ԣ�L��Wjh���S�#{lu����ت6�el�V�����>��������!�ū��;�(����?�K/����:8������byi��A�>}R-��fK��UY�F�_��ω%]����U����Y(u�,��[��{�������*�M�=9^E��9۝�m�dO��{S�{_����wlS �%E9(|��v��I���0��K?TH���[׮h����9���I�ՕEloV1PƁ�1qA+�V����/�h.�rXZY�b�&�	t�^���=/aeBA�5IP��ફ�7�)�Ue��S�gO�;r2�3�NC��t��1]�	xN���8f�G�3��j�vs7�]�V�&.wF���b��=�Z��nk[�����_�)&ff0*`��ɣx�3O���x�?���|���q��8~�F���%�`� 0�9��@[b9���	����x|��A��t� V/�a���2������fG�2!��Qӥ�M��(��X���I�igq�憌�*�0Y�a|��O=����%��7Lɫ $	
����î�� e+�� �"s�5����ͶK�4;�n�@�+�dl����8�����~�����,���_��"M���ͽ
n~�-�[~9>��	�H'��M+�
)~zZْ"U)h`vbO<0�J��+.㵗��z�{�yLLM
�u�FC�`uI&ي��C���I9����ymmq��	��E�s�<q�nFCc�4kU3��s�A/�D�X�)-LO��~�� ��zi�t�ZU&R�(�<P,���Ym�6�9��E�:~ ��9�����._īo������f2�:t�="V�Xr}1VL�*�o�bhm\���g�C��9" �4���p�y�͌ㅗ�����H����+א+MaC����'+�����3h4Ž�����O����q<��q�M:�^�������:������������>������_xG�C77����5��ŗq��-\���W���W6�_|���Z$_F���l�Ҡ`t[�\I�)�FL�T-#֝��3g�\;2�9WOlNإPd_�M�����$�-t�"�=Qn��qr%a����Ɏ�װc��W}l��G'�z/`����{�����=�r�s�'��A8�����W`���:o�K0e��Դ��L��bs=q��Y��vv�@�$y�@[�~� VYq�1�{|��H��"��?��ݗj;�68*~.z������]6�)9�ږHy��h,{]C��<���l�sr<�[o��X[���8x�j6�o���!�Ԫb�eqpb���`j8�텋�s㲸�8(�3=5���8���XYŲ~��\�o*e���	���އX^��'\���ߣ3%�ySAJ�=�����E��M�B�����>_�\*��oٓs��Eon!6qxrJ ��;��}��,)�Jx��G��O�����ׄI,J`������E\�|o���6���7�H���9s���cC|��wp��%�'�kU�To�駏�`�YkqaCS'��Ņ�Ǒӏc��e����%�bmߑ�4W�������(���΋��7��`���3��y��?�Sԫ�=-��rm;����'���~f��bIOctrK��ÖszQ�0��4(�J�-�j�: �15,4-`�A���l�ru]�й��D7u�U^��V����$�_�H��m֣�{˂�����Ж��g�j���U��l��y;�m�*��y��j��a]�U)r���_g@.�2���IpS6�[ߨ�鈄f̌�k���[r&�t��14��������/��AJ[�DM�L��g���-�������s��ik͛J+�Rim��s�u�a��~$�drdӰ�hl��o�H*�V���&�q��8��b�����.fe��(q�ƼN�r!�¾�`��"&h� M:��cJ���CGL}����U�����;U���4�*�L��2��~��_�Cϕ$`��X���2��3M.��&:�m�9��a�B>���Q����8���:�<�������C�22jKD���s�j?I��N���^~�e\�zo�����q\���K��?�k�ϟ��'x��1	�䥿��Ĕ���jq�<0w'~K�al���0v���dlB��ϊ{Z��YT���attL�t}u5�'�n(��5R;��nV��9��I��0e�S��A/^�����-#�[V���d��(��A��O�&�:خ���@�W�Ϥ��&,��Qd7 ��[F;?�mz���ܯ�����ݡ����Et��&>r/M�p��},+Fw� ������9�d�?���
L�o�t44év�K4�Ѣ�Ѫ����g�zrV#!yN�=@��&�o�o�<��5lM`��6�n�k2~��a^a�CURs�MZ��}8B?q{l�y�M+�����P���+�LG+����{�M��T�(�S�bdM�8`����p�͖�2�(4��,����HgN>�'��굛b�a���ҀZ���e�[*� .z�.`&���~�y�/o��w��8�CX�6׵�{Q�� ��v/LYg:eVM3����[51_'UZ�L-Om��z|x�z���3G1R)i��7_{��!|�뿮���I5�a�~n��K"ˑ��=�Z�|o��Cj����K
�o�����C�U���7�7x��ַqQ\|�G��x�Ӓ�L��C2��c��}<vB'0�A�V��֢��X�a+���$�Ʀ�!�������^�����>�ڣ����,NT��b�$����R�ƚdW:K���=�2���Ą;�zZϿ�����|Y�M9��1S�\��o2�}$;a@�v%�軀�0&	m�@1TA�>�r�d�H���B�`����Z�S�u��EQ�� kN,/�����9_+	i�tB��i��E[�|�w{�@Ğ��D�ȩJi�
8m�h�7֟��i+D]�#qw�p����f�2a�P�t�a6a�}�-aϔ�3)�v�N"�%�<�e���qw@JO����5� �t��H���ٛ�$ J:R����;w0:2�U@�kj���h�.� YK&O�֝�hj��<X���88q/���y�0��c+��*0u�X
6m%�4��\3j�B����P҅M&:�>22��*Eq�+�ˤ����oᡇ��׿�u�y�!1�+�jRFNe��<R;bNɛ�� t�>�����W��-9^~��;����NN����9��pE�KW�"#����A�*�d!��z��|oS,WZ�Iݢ�jh�A��6jm�S�ͮ Y�����.6�j����wSƟ�c/�F����}�8A���z������7M�xAM���a�=G���{��9'߻�0>����hbR���d��2)��02c�I)U	 �9�m�vN�0�/ݤ��[I��-����.���g�`�����8����h;����:5��!񞃴���e\�$6+���d�Q�����8�
x~�#�ϑ�@��s�rp/eʛ�!�m1�Z��4��H[�zD��-��y�Y��Fx������6�M�p||sss����)�	���E�+C#����3)i"�o���g�T6Q����nyi��,r�E�� �I���&677t�TP�ͳ�q彖�<��D�j�D���<nW��+ixx/#����L�j�����m�V �U|�FTO�^K������ (�)����/��C�N���o��GK�= �Tָ>v��� �
�D�3].8){�|�7�	���q|���ť��q��1�p{aEk�3�2&eU�����S�[��
�\S�%���)}���8���d���Qȡ#�@[��I�\)'Vp�VG�,�恞PM�P�����9a� W>0�-A�Qqr�7�͛���܃lF,ܮ�a����uY8�~����3L
Z���˘�D�Td��.d4#��,rw�Y_�%\R/�����K�a�->������]�{x�z�ز񬗥ߴ��
��?	%n�-��Ј��t60c���y��w\_���%*��Q8H���8�5"BM��иd~�vW����g�H/�LK�Z�֐Ѽ��AF�������{Kk�O�*�u���TF026�\��$*3��u3�����w,~�t��
�֜�ȁ��V�Mrɚ�1l\��m��Tʪx�y��J�d�uʛѱ��A`V� �%@�X��dn��)��C��U��E}�������)��^C1�äX��4Z]����8rh��~�<��aW�0rgv{Iԁ��'W�߸L�}�����H�m��9�-�+�}6��kh4[Z�Z����mx�1����d^Z��yl�*�.erF���y|U�g_&��56�ͫ��ϵ�骚W뿣߁$��ۤ��gie��Y4�N�y���UN� �@a'���
��v�'�Q��&k2k��N�t�wLr���8���u�H���7�r9�%�?'Y��\�~��?S|i����|�vn����)�Қ�ۿp��L���?o
 ��E���U��-���A沾z�î+h��9{��u	5�@�-Qo�&d��\��]��<Y�j��e=����#'�� {��JsL?Z\5��5{�ɶ���<��17���3���3�{�$5,RQ�y�M-Rv�Tw�z�2д�8vL�0Y1k��k�u���IIK4���L���S|�Vi�[�����C�T*���ju#����b��~�������Z��ăm2B���.�F06TPP�u�&F����7��<��|p�:/���Ν�%�r���Y��s&xo~-����O�����~O�z�4b���xCk�~]�p
YU���K��hiC>>��y�����Z�=�(y
��׍ܫ�Jv�~kV-�F��S�Kg,�8������@sg��D�}�F�/�OG�G��cO᝷������F�&�.�c�[{a٧�w��3)(.�Mm���-�5�i'��Ը�;�ҍD5.��#t�cſ��a��)u�2��)��� ��4+�wF	7����L&Y�z����Qx�,gޙ��f'ش�S�Q�:��k6���٨�0M&�u�]hAK�5td�`aߔ��(h��h-���y���#�:\���֖�h2��E*�1���^���=�=�3���,��A6����9�J<v��S)|�-��}���@�h���Г��5Ԕ/V�Д���v�N?�	q�뭚&:j�C��*��L�uC��)P�0��nȀgq��C�z��k�F�Sw�Vcq��vꊕ:48(7��� ��Y�eۄ���nb8�B��r������e&�Ҹp����+_�g������Fkl�裬4fL��������T����������
2oV�J�gs�c��%ۡ��n�����d�D�.^��B�)���؁Z���p��Z�jݐ�Go�Z���{�R+�FcX�
���=��	�2�����"$ѵB�տ�������^��*^E�WmX�X�X7.c.d߸��Z���_��=�>iQ�"����:��&K6$l�� 0�ĝb#^�3�N7��:ˬeĽD� v��J&��w_��%E��<��dBɝ�Z�6l��gm'���s���i����"��2<�"�L��\)�S.�`�����U��s���K���+kR�/*cc����xJ�p��n޹�\�����ዿ�y�>qBiNCb�1'�U��`�.�cmc��� R��*=���	6R?�ƱͿ;Ν��5����8G]&ɦ<���&gby}�K���`���5A䴽M&;�6�+ώ�icu1������z�2����
���iuԵd�\("�ɍ���Շ#�~�G	
�lRk��\��X���,FŊ���=83�O����P�%��R^�w.��ی����8N="+�yY}����P���2�Q�J�5X�d�c�&���^�
�L�$�k"�`�s}�M��&g|�v1� Z�h�EV�O�u�:�Τ�ɡ��k��d�=�����z�����Y��ZYu$+ޭ���s�F�>!�=���Ga��da�젣D9zO�1�.�"�mb�Yp��eܬ�։޵��}�(�:�&B�|���6B�(@k,ι�.j�&	���p�O����<o�}���dH��X��}�-&���<�6���|����H�������W��,R9o]<�s�Vo�X�d����>C�gԕ�S�{�R���:~��kx��y��v||bR��~�{���ϙd��7��?�t[���)��c=�݁�xN}����iD��N#j��
�GUz�y.7�*�xke��<���_�����2xS���Q`k7�u¤�]�2�v&3�t'x xn�԰�Y��v[��rJ}qط��a����nC
^��=@�t5��\Sy��T��ᲾXO��3�S�SJ*l�.�Ϊ��؃��ؑ9ܹ#��nb\����A���;(7��`�h�0��������r�� ��F?[�վ���C�9[0��!
_<��X��<6Wxz]��T��n���b9��c05;� �Q�-����+m󼨒&i]���/s�u%6{�*~�ן�{%�YP	B>t��D���,�7��)IΛ8�$�v�d�ĻalI��E���dZ�ݝ���z��~Ԕ�a��Vm�ڕ�x��W���� �p��f48j�3,T�${Ϙ �5۳1M���P&��&�s��{�����ǟ���8�����Қ}�P��#�����HC��O�'�}�z_�7�5u����\`�xk^�<���!�9���*�~�}��fp`zŬo�������0�V�p]�תب����ĭ;�b�r��U݈O�+�Y�Fk�ܓZ;�m��ZPf:�C�Q�8�1<8��BW�%���g�X�g��ݙ�D�c�g�]2=5�C�3�_X���N=p/���J���^�s�l9uH]�U'��ȝ���Ye.g�F��qܳo��[�	��c:���6Zu�,�ͧ����m�N�4�
�nT74&�37���A���<�XEI!D �t���2����}��b�M�_�UN~��Ԧk]�[0���Ҷ��@sz��v�ov��l"���" �?��~��<ۀ�=���9א0�����0������fB8��Q`zf'O�V���G�G��TK��"��pYn=^���ѵ�H�-pDWVV1����C8������Pj�f�.�� ��c�\��"�4�;�P���mH��[�c��n{Y����@��?uM�Z�i���xYV�\����<��S��l����+��v����v�3�=�*���
m,��am�*�0�>��z77��& B�S���Y�s)�9�?=����0j���
����I`��V#�
�`3I@N��N��xH&\Vך����a�@4�?��7�x�sY:0#ܚv�;0��@�ڶƧ
V<��;��o�������T��ڽ�f����E"z~u X=b�@'/]|�H�N��K���<z�i�G�C�O�� ��#eNYM��X��=H�Id��c�_��y�Z�Z �@�a��S\z�xu�D9)�O/1�v݅�`w���_��=j�w}kU�`?pZ}��1*���T��M��C���ᘌ��ps���8��*��W1(���_Y�6�=+*۱a�U�f�t��]��ťe� -�:���X���wR])W����B���rekY}~�����=�������G�,��U� O�XBGܹ��*.�hj���3��*r%\>w^\�ױtg����ԘX����Q��07�l����h�{���)���Lؼ��@��i�q|0�ͦ*�;2q�&yQhSO4e\W^��Rf�ewO0�N7�ر�� ���ڵ�y�ЂO�Iz����1���k�����Ӹp�����F}ϨU�Re<gB9�L����`�s�LZ�{��gt]�m�ω�h�JE���_��+���������䐺s�$9I�IEx�6e�fSm�����mk�k��B��;���c茻��~w@�%�t�z��}�I�t���|xw;����0a7yo�h�w�A�^#-�����`�RZ���xu��<._��9^;q���m�
��u�D�����dCpl?NZ;Ɏ��ctl�p��};�>*`Z�I��%��K�����N!?`��K���Z�]�{��B��Kaf\[]��BA��d�YY�;h�=�g���O�����Ν��x���'�k�� ���T��`��v�n����#��2�2��;l��Q�94�El�����qSr�r����՟ �Z�NC3�#��0�h�|�2�g�0�!>9��>tT�����[uD��Z��ɭ��7�㡷����f�y�:bg?ᄪu��><���֣��k�rn���1>}
o�u	��_����(*�5۴RRJ�c���I�ef���Th�L1�� ���ݝ:�x�I���M������7QڨqCKuq�)�pS���L�����W��m��'t����gֆL��޹/G��W]|3Ҋy�q�����Q�@��\h-�)���7���7o�ciiEƦ��M�"JU�5EN�o5����hV�-㡤)�j5=9�eq�G�'��x�O|Hp�^�2%�	������y|��e<|���>���?���7	�&ٔAD`U	4++G ���ۋX_���U����A1����֭���O_�_��3��y�1Y������&�x	W�;�b9"��s�*4M�2���hZ2�+@�?Pn@̃����B�U$h�s�r��%�I�D)=9L�ɸ���KiKg1�U����y�{�)�T�X�$�H��dx&v��k?�\w�Xv�Fk�B�;]��*�y]խ:�N<�n^x���+�I�8!ו\`^_��B^��.Ҡ�H��?��{��d�����_,؇1�kY�k�k���v�jH��6��0�i`,�TJ����v��.45��w�c��>:��5���k�v}�ZTh��SC�QT��nD�J��{����OKё�I�g!GK��|���V�p��E�aҵז�r>,k(���1Т��/y�|_-��-o�0)��※�p����nQN�X�۵&>"��cqy-qeF�y�xq��Q�d ��P��m�"�3���M(��@v��ސX�-��{g/.၃q��q�N`�X#i�כhĹ����~�4z9�B��Pm���H��F�W�:���1Ԕ@5I�d�$g�ڴåO�4Ѡe������;��r����$g���AME��*�����梓<d�7".���<�=�llbe}����#Z��R||���5I���xHR����3��\�75@�v!��BB�3�y� \q�~'�U�3�~��VB|��ϣ$�c}���K3O�z�-9~'P�Rf�����H0?�kQ�2�ɞ���"ի����8
b�,	2fP�H�d��4����b򔹈{~/:. i,b[���+�Ϻ�I���꽱8�>�;s^~W�����ϖP�xN�1ci8�1M��2����頝q��7cC����F�bIH�f��������H���w;*��2	E`-KC�i�� �=p╖�ꨌ���ӖWC��1�R��%�o�>��`�cS�.r^� 1I���Sa�j��V���+��|�R�ř'���;U�ݯ����1?5�t)��69i�t3��r��,�蛕���d�	�t�z�u������J�Ә�M��F�����R)ib�3�n��L��4t��[�4B��51�������Y^��p�<�my�B?� ���z���v �a* MSBg������E��v歜x��������k7��U�" P�֗k(Oߕ��;���5��g͹��ޣ�W�;�
G����'�9i:@vkDm�̽��<�W�hh�?)��\vg�[�؎���zTv��e�܂Дj��eWK�z$�z�TL�o뻙���rTm�'7zk�Pu��^�~�W�a����ˋ�.���`K�LV 8tG��B�K�.+Wtp����u��pQ�O?���9��{x�bPZ6��b	I�@����Ɩ��Ј�{�M�,p�ڤ����R�PU��VR���Ϣ�N�=#�+�xFǒ��z�ba-n�!S�"7X�ϋ���(��$�,od[�к����]�@�}�_Mh�3��J�I WP��!e�/<>+B�c��n�q���ʡ��Ĉ_�K��f�IPNG�!-v1���vK].S�ohXᮇź�����#^��]�Zy���=� ;�K�8�+�����(Ǆ��ܾ�������b��x��'ɼ�LZ}I`���:�Hc}�r�%G+�-��.�;��!��s���b\�[�XF! �M��'��?oֳ�IFy��rmu-qo�����9W=�,�$�we�P�8-��T*aE����eL�@E�Ye48�Jf��[�ذ.�!�cǏctbJ�Қ.�[[[�y�E�x'k���d�����5VV����`ڦ`��c ��i�T��ѣW�SlR*г�9���qO��4��T.��l�8�;���]W_6�H�d�
L�Wd�E e�&*P*���� ��j��|4h��i�̇��F�U�qͦ�k(�.o.7Qw�'��y���<�	�����-�������yrϱK	kQ:����g���,2'R�j�DV�ݏ�H(ݨ��Kĸ�E�M'w��QYa*�:���Q=����nTaA�x,�j�x1�_���l�����n/NjPՉ���\r�0yv�v�OB�֒�M�E�Ac�.��r���B�D�J���������2�y�]~���s�O�2�Ź���~cG����(��.|�����	��v��P����y�ˋa�q�G�F�b^\XT^�Y3�\�<�h�5�����j�5��=|����fS �S��`�3�gr����XF&���2�V��/S$�
(d(����k�f8�(�4t��!l�Ĩx���s����&��<��xXo2�Ӳ֜ig�8���j|�ޤP�|PίG]R.�<)%^�@�����ԏk���L0ϔڕ{u}]cD��$��P�hB8�܄_�(Uocf=��*��T�w�	�G}Ë�\���Ŧ�f��I)5$,4��p��%V0���5��LKՕ�Z@O�Q�=C�j�A������9Ľ@؆��hv[��{���~b�a]�j�WEc�.�3ܻ�#N�l��7�S�	���S�F��s*gY7��$�`bjg�_���%�iLM�`P@�#$�onW1RƱcǰ����^��)�NNNbE�f>獆��ٜ�v#�BiȌ��x��me�[�~�e݌�C�Tk)���N���Ӟ�Q�_�ڊ<�M��<��J��>��=�⤀R�S��+�ժ�0�k+�_�w�#�,%��P+��0�����i��l�R��W�qE�b��9+ �xUƺ���Ygt�����"5̐1ۺ |�[�XHCٴ�{�b���pMa��L�4v����n��/��f����i,�]F{����Ưh\�I)��9�6�2��dJ��G���ыJ5�J���]�N�k�
K���z�{�D����2�Z�ւ�@+L4��/���Y��[�ȳ��]�B�hy.����{fQ�]�$/2���k�}Nh�x)c�2�T,�����ￇ�9|����SGPTwsQ�p] �r�<�*5UkX�Xǵkו��v�333�p�<Ξ=���Q|�g12:��v��$��kG�T*�0����'(y~�UKD�(��	Ž�n��[U��[��~��T&f�+���m��Ԇ�N�&oc8��TkOJP��fp���µѮ�!��T�&t�	'#�GKn^�'^�Y�<j�t�4*�A��[^^1�Y��Z���h��5>i0u�6��5y�jX^_S�.NiCA�����BMԹ��@�P�{��(�t����$��O&�ێd�;e����֪��^���5:m�:͡Q��~;kۚ�
�^������w���1���gϤZbu�/�����y�Q����Ş�YH|��RS��!�b'w�8���H�$q\U�K� �b)SDS��z�
�ObhxH%-��d(nB,K�t�J�ɝ��ړ�-�>�w0<4���d,��UT���b��Ʀ�\'f2�V��d�=��7�#�ܘ'nq}�ڦ��ۛ��[Hy6㊛����q��,3�k~���q��E��YqZϒ�����(�<LT�\�&A�_�m	kG�t�ʤ�Qy��ö����`cuE�kyec�b�Z��s#
�&6���ǄR7�B�F��������d,����he��n�L��i/���ؼ�\;��؂�w���k�ߏ�gg�����C���{�T��3� e�bO��w��±> �~�}���j�����Go�߹��g�ݰ�x^��Eڰ�!��iC(��>�3�^Ԫe�f�́�[�܇={�΀QQuT	z��i�!'���ir� W2M�6�7�% �8���Ż[���
�\��a��
j�m���kwM�o�������]][��n3�t_x��=�2�|�oצi�I��
J�<�Aq굚X�u-d_y�\��b46R�9!I���0T�ڽ�����t��Ƶ1|G�����#�[x��S�=���3����W�}0Z��.ǯ
`5Ik��)`��m\�yK{*Ur���L�)���Ż�=F����7kU�YZF������C)�U�fr+��I��8b�&�=��f��8��LV��e����H��
�N�1"��|���xu��F#�f��31�z�������uu9�^������g�y�Z�gDq��w�=�Θ6���3�ؓ�.߅L�4��v¸o�����&�ͭ0��	vc�%1�9�r���'����
��H�16OII���>��c���b$%M֎����E��gk vz��U����5Ň�
��p�;vld)�ſ�J)�Rl��������n
�頉^uF
��/<�SB��U�4��UA�7D)��r�c��W��'V� ^]����U���4��^�F��t��*%��z.�dH��f�"��iq�kߖשּׁ���K����..�ܝucRJ)���o���������t��c����~��u\�qA6�M�ב�\A�XhFC2��H�,�)m�'p�jSK	먿�z�U��*vT�c�iY�al��v�������0q{�(���p�G��,�$��K��U�?�Z�{w�C�v����{�ek)]���1�u�;�i��Z ��c��oɏ\��'�	���X��|V���X�[J[��������|����kJ�,��hI����-ܹsG�cc#�^}eyI޻m;]�������rԣ��F�U���Nf����5Oɦ@�p�.�T/����y�pqQ'���h����G-(���]��_����!���ߡ�W:�+h��A�F<wt��j3�ʬJy�m�.�0�˫XX����4F&;X�}^��ѱ1L��a�{�fVh�}���Y�֗���������>67�;��@N\*/��k�Ώ��h@J��N��Ϡì�(Y�}��)vi�h�,8�Ne�U7�-��t����0�՝�]����Oү���{;@i�m3�%xq�E���-'�������u��.׆�����߽�7~^���m��D>�+�����ʐZ�;-a-��uqѮ�~Z��^��H[��ban�'p��Q*�p��u?����e�6C�0��!!_�
Q2�ڔ������Q׳-f}错���÷噌��F|̌��M�\�wj��V�d5HTw��)�?�7�w�&�kv���G�\�9�Z����!�5��� iO��iq驙|�֢v�F�����%\�qS�*Х�S��|"wW�{�K���[�:��Z�����˘�r�XZժ����*������-�%��>���s�d��a���)&?8��f\|�mx�\�{��e�w� �ο�'������;����{�(��w�{6\`���v��w�]GD��ݰ_U^�E�ǎE��N�6Yv��DS��ɦ�N���41#����ݒ�[]��<--������BY5)V�K�U�����zb5	��b�p�)h��s����j��K�)��k��eQ�yh�v���9*I��$ӹ22���l$ѕ4ߝ�ꬽ��(�D��Ce�Ω.�k�������Q��[�t�sRgs�eĽ��������a��a,޼�.^��� ��1��J��Q0f��ml�w��m\�WK��+7oʩ�044!�g�Q�Z���Q�<�1��]'v���_{K,| �	�Z83�%�џwk/\H^��\�=O�>\�����OtK,A[�N`$"��Y�	zZ�%�um�`g;a7���بw?[ ��7�9��2��I�ػ����!jY�l��ٚMUx*����h�$e��� �Ūe��z���7o`qqA��߃`c����[��=��I��N�㪾m���Oզ@�sh����j�W�\�(���̢���Z����%с��i�kM�Jc�6Қ94[�*#�5����h�����o�ş��Ƀs������k�I����	���7{M,���}=p#SX_������M<4{@���O�y�<|߻���;�t��K�+x�}�4���9�\�WZ���$�̀������E>�i��$	I�l���Oя�w�<	��22�mH$iX&�Ͻ� �K�g' ���u��`���cA	��M?�,u5	͂+���|g����K��?�)Ƌ���{���$c�ч#��%ͽ`�W(s���pe��k⒯��4��P��2�L���?LeU�]׹Mu�i�~88XV ^���^�0��E�L\�L�A��Ǝ���$�1;7Қ���L	������a��?�����(�j꼫\R�V�0$O�3�_���Y�GtׄH܁�Z(L���MUe<���]O�ڇ��`\�m��鲳gL:5*7\,��7124���
�N��獄� �Ⴧ��-lͻ�&�����j��.�\��pQ��7�}k��� 6�!d�?�{n�$�/�M.�^���4��Q�OɸWb
E�ƾ4H����I��gubC/���L];�X��Ϛ���K���3ْ	/J�щ�������_k��a�'.-:��|�s��qzɘ{��}�0����i���E��Ћ��y5ʚ�����|�CY��1ʍ���1w`[B�ju[>�G>S@K�]V`�|1��Ō�kXX,�1=>�s鎀�Ƈ��5L���D���m�)7߂+���S��
�[��i��W�c��ae}be�����{�u嵕#�FQ!��w��l�[���{��=-��b���PÓ�n�|/W09{ㅲj ��Og��n���zm�ڭ��t�I�
bg� wS#���|���zu��G�UuX���Y�5vo��/7�K7n���kה�A�����˱R��4��mƈ�FZd�!��D�_�V��:�g������C��:	-�G�ш��!��@��� ��xv���A���' ���{�c��~��^ɦ�z��ߏK��]�k��K�����^��Ѭfo�X:�6 ��苩�}����dv�>��h�6c���@i@���9��|���|nb|)�t>�Ρ�^+���i͙���6�_���ј(ۜ3�?����;Kj�RI��-R&��%�����L��hq�_��-ȵ�*�[w�$��x����e��ڲRe�ղ>S��&�y��:m�
�V�f�Z�C��\�NG7�}�kh<����*��@���e�\XXR���Ki*�*0��S9Omi�+3W�|���y?5p�s'��l��,���h�p��Q�SI�mz�#��=�ᮟ�0�D���_ݕ��q�k/��(يYF����$/�C�����? l�T��%^�����\�������y	�ܝ��鮻�o^.����~|~L���_һ�o���)�/Z�њϷ��|O^��F�B��*s'�(�	�V��{�?p���x`�8�Ъ�#�a(I�M65&p;w��57�>�M�������(�Bʏ�+�Nn��m��V���1�J�1oz�&7�Z+J��:�
T�8���lNDt�;B0�{�q���K�����Fb#Db��#����A����J��)&^����k>aEC�l�n�F��ڡ�l����J��xDc^�h���J�;)ݚ�-�MW�lz|��>���إ�.K:[,i�}��{�Ա׸�W4��6N��e�uhϚ��!�������Of�V4[��BMi�p��rMi+EFZ'�M�ԅ����]p<Pdo�О���䋆l;�L����I1#a��xM3X�xKާKv3��%�\��AzR�M�dR�Aޥ
��C�jӜ^L�T}���X�����+ZϮ��_���=��>{���&cʇ��{
:+��~�vhU<����)[�����.xJ�W�9�{��x�Vi�M�����
yI���ԭ���C�,�o�pɧ�;�	+w�5���r���9��^n�<߮���H�U�|�-m��:�KiTL �h������x��I��R�9@�Ye�Ge��21
}�d�C�9ʏ���c�
�8%���]f��$^��MK<���oZ�ݭ����|�<���fRX}��O��ՄD���b?
�S��۶*	����GK8(�|Boo����.�laΦ4�4��5k3���������
[�+��B|�8�SC#:��KZ��=?��w3J't����קlĜ������zE�?8�'�w�l�:�Ԇ@gc���[!�Ci�K�hOU�ڣh-�7��4�S��t�:t+�~������@�d�J��
�d�dТ$��2�	H�Oc5(���qV���X�"��u1ߩXp�d^]���e����_�Kz�Boz}A��?��?�-����Y�N����Χ4�4��Z��X=�Pa��R> �A���s*�>�<s^`7�B�}zEgW+�~��w:�5z��2Y��rM���������{KȺS��3%o��F�ʤ�"��l�$!Ҷ�<'�,s%(B�"�<������~r��0� ��T�������*q�q6���,숻q:WO�`T�X+��DZ�	Jn�~�k�S�'!W���iۈ��KŃ��kB;���b����N�u떽Uj"�EI0��p����%��i[?VKZY��·#u��A���Ns�7�(2#���!�	�G1h�f]�?�}�^�+:}���[}���vm�
g(��u�����IH��	s�%�Ő-U����K�EǏgW��{�=>8���B~��{B 9e��Iʘ��G�V���H�!?�qJ����dE��J� (ul�IV>gwF�DjO�w=���2¿#�g+5j]k5x-�M&$e��8ea��k(	�Qi� �Z��-�X(�����r�/D�P��E���z��o�z��O��Θ��<�-^-�i��ӋS�C�A�Ȧ�Xz��(�t��BE������ؠ��(�$tН�&51�,2��d�Y��.���`nm��bÀ��q���a�;n <�J�r\m�k�����u�}}v��v��آt���z���0�?qI��$\����~g>h��	Sf�	M�ͧ�r��1KCвX���T^0A(�M���J�$~��#�b���Z�(���+��[��*���ݧ�)�lJ��CfaL:7[L�F�R�,X�����G�_���y�xc��_��+�ݛ18 �D�w��[��Y�,����00J�v�=v�k���`_���r�9�x͡jg{�>�-�ƒrI� ��`�@"ܢS��>�g���Ԕs��oO��� gO	+�j�J�qpٸ̭z��$��$��"E�o���5��ַ�6��w:��Ů����"P�J���=�]�(: i����gT��t||A�o^�[�G��%���v�u;N��#K-D#>桕@���-V+:�^���M%S���"��q1	q���h;T�.j��H�ܑ�����V�r1�y
8��:�3��W)��n�H���R(��S�BP��)������u��X��Bj��Q�Ѭ�4���t�5�5.
W勵�F]D+tn.B7u�@"${#��g_o#��6�	��58H���]_�"(��$$!
ػ���ХN�Z=����W����,N_��P��B�I� �d�4^a��P��.��uu#�d<猍��$asg�6|ԒRQ#j�	W�m��΄�R*dRQ�$��eZ���@����X �I�?�x����3������!�Q
�{�w�{n���5-��[Η���h�p��"q�l�|�<�����>%���������z�@�y<u�U�9�������%,��'s�p>��Xm����"L#uAS�4qUHL'�M���� ����j�Ja���d2����^�J��Y�%O��?��-�0}5I�����K���"����|�oJiV@]*��Ӯ���NP7⭴�,�F��"�'d!D��C�C$�Y�i���L`	X4o�ι�f\]Y$���n�G�h,k��H���N%��:��X�y��0���%�lC��ɢ�l{�=�)d
�z�5��Y�斕��xX�^pm��4���0_��8�8�y���☽�2��R�8�)�x漵��k�P�k2,N�ɦV����[�\R[Ip^�)�G#��T�`�����43�s�Ǵ�eU����� 6<,�ĕ,JL�Kf]˓T��<��������������;��?��Q��
��,�y�l=�k^��Q5����Z�_)�z��FO�ho��B=>�y��9��u�x���?��;]��t�V<ApȀ��p^<9�_��b)��rB��,Z6�d]���s��Tcu�Q�z����
�K���_.�����X@�8�x�+~��ĺp@������&�+�U�EV�Y��|�=^|֬�S����6�L�.��Cbh��w t�(@--0F��H_\�eeŮqk����j$���f���׃�5ĝ�0ۀ��1���}��pA�J}�(���S�=�de7��;����%?���ab o��ӧOU���CH?ذx�z��:�:hU%�pC�1������|�� �5���c����,D�����%�dY/K��Y9�7�s���v�7Jo�8`�(�� �}���x/�b�%cp~s�ct(�$�����|�B��5�b���\��;![f�F�5:��+��P�$�&�ڬ�n��A���,A���Wv��s��6�u�����yB�zE{l��Z^W'�?�9�����f>��2��V������^Nw�`�w��W��k��i�t)Q��pO�R�H�UCG�=�e�<�!�X��_���k�5�޾��`�n�gtI��t$�5m��z&��(���7d���<G�|��цg��%�̥p�t�)���Zk�t!C#�f���1�q�i�A��%�"���־����K}ȋ��s|9����
��4���1�(���9N�1ڜ�c�@lZ��|�zS�V�v�pAI�0�r����CKx^ ]����	TX�6�ִ{A���1�0r��ҡb��[0aaܔE�]xkI=g�
��s�K�u�ڗ�ٹ��^��ժW��R*4Κy�&���K�J�4>�,h��k �����m��Ƶ+)���.{�VcXyU���Ƭ�$qy�q�Ϡ?1������R�jL ���P�4oI��(3DF��<��RP��_�?n��i���_���з����g�Yd|X�H>A��*���uG FAn�͂j��ݭ}��{C���\|��L����l',C��{N�S�vQ�8
A�߷~nT98a��N ��Pr������@,Gs�h]��d1�"��J��P���A���LF8A8���H<�$�;��rN��a(Va#@��+r���\S �潒/J6'���A�v�w~�_��X	I> ���/;�{���-�C�cH�sI4��RK�¯=�WlZ���!%�e%	�!l�*���ז���pҖʭ-P�8���3w5Fa�\dFX#`�'f�̄�q���{��"w��q��j���VBν֓�>����ɀ�;2�c��$P�v�X�x�L�[��pP�-s'�cR*����l6C�(QPP4y�]J�Q�lb7��`���kV��R����و�ޣ㿒�5_$��f    IEND�B`�PK   �F]Yo�>��q  �q  /   images/2cd737db-51bc-41eb-8762-f3273c40eae5.png =@¿�PNG

   IHDR   d   �   J���   	pHYs  �X  �X{�M   tEXtSoftware ezgif.com�óX   5tEXtComment Converted with ezgif.com SVG to PNG converter,)�#  qIDATx���d�u�+wuu���9�LO�   $ DҴ��l�Ғ�//�����o˖,��%�f	H�� #@�<��9��t��s.�}^������*LWx�{O>��+�/�xF�`�5Ci��� ��ɂpE����0�(M� ~>�ؼ�Ϡ��E�h�slyh�lz�k�.����ޏa~?.�7*f$c躴W���8��F����kX'L�{�������������;��|O�ԏ�G��Iy�7�r��f�l�)��ϔ��_��R��zmU���˶ғgsy��YX�&ē�Af\|�j��,������XC�����B����c����
�k߅��,�๸zb$?wD|roS�r�$��%����׭�u���fHL��e>��0�w����q�W'3�����/��'�A�s&)+c1fL�0�y�����xP1�O�^j���-�^�^�1C�ɰ�q���K�pq�mȘ��r�H�z�Ɉ�3��e�:��U/��_R�|U�J��g?ٿT/a�}��=�^�׻�U��;��ں��>����Q8Jl�%���3����9�}`4
�JSN��蜼a&���~���� �qj5Rg𚚘�"dN���T���yo�x@�K�m��~u�fܱ��F�շ��jZj2��.M}�W̐{|���O�aځ��]?����m���w��+������돖s$f�݊P]����=����A�g䷅�Иn/1���V�O��߁�����͙MbN'(ok]g�V!.��%�7���PO99vje��M娭.��T&��&����1_XM��T&�Z�u7��²����Ȍ<��;]�/�^��_��n���y[gF��~��a��g�`�u,�!$��8��b��� �V3b���J�*��ho��4�W��^Ĥ'R ���4�Z�X�U�V�nW9��¸��]�82�dL��Ɂ2G	l6�.�z�Q��.��'W���D0���w�_B���������m��� oc�$�}B'�{��[�j��>���7�N����oe{�!(ťQ��/m�+a�P8_(
���:~9�O����5ÙV�հ�5msAL��KHnv�Q��t�l�� ��UR��1��.�t�Ӭt��V��`8F{U%&� CA_�41,c�g���/�h��"�X��AӮ���E���A%��"�_S>�&u8���ΐ{�k�z�q���i�����-�f�ɑIܮd�_�qkj]��d����"FYi)�������I��9,-�J�8�N�J&10�E8�+��E�(ä���9�X�xnIf�[�a�K����+aK�`���]�h/c:C��L[ZfDf|S�6/�.�������'S��T��<"Ay�����>̏#�b^¼���7C�PL##����`�8�ל�L)�a��d�d��yJV9�������p����_������H0Z�����[�������Zh4/�x�������TF�\r��p�e��lƺ:7�?�+�I=�'��=WE4����ai)�^�xj��e��D2�٫a��ӞP�?>'
��M,a8��A�#�Jǐ�]��8����A�uU��K����ك!�?�(�[��,8�+��8�N��[���Ħ�e�+�2��,��U�eQ�>y�,�͍5x��E�è0����@�W���U.~|c���*�Q���:�M�R^���"C2�)dm�I`6�5Q8��=~�vZ�J�a��#�?�}.4��3i��
Z� ��hi־>Z�E�9�ECi���9�F�/d�k!Ys1�a(� �l�P�L��T\-5�ƹ(��4*��̱83�3?���4e��$�:sB&�@ځ��2�sFe�L��,N�"ڮ�Z�I�.���nRք��8�a��	dсH%����Vem��]�z��M81<Y�3�$���i~���	���xlp>eyݿ���	*��u@�o-��S�#�P����U����ؤO�0���2Md�PVQU}7��~ e�b��Rq\<�.�~S��ȴs�V��*$��]��OO]Ƒ�qaC�5e�p�,�V�,�A3}�@>.ǂ�妭��ýsT�0S���3^�8�������Ճ7.�''/#O�t�.���!l�p#�l�[Mv-ҞLFP���>��z�S+�S�Ȑ�Qgv��(�6�:@���ذ�$�a\�tX�y��'����E�ꮀ�j��3.���|D�������[�aH����7:E� =�DzQ_��1b�9�ڱ�DF�X�8^�Ua��nU�e�HT_ ��U,c^�����(�����dZ9�a�[6���5X��~d2i���V�l��]"�↨�Dj��S�+�4�n�����_�4��f����m];p��	�	t�&#qE����كjFT�m����;wh��xbY��E��*Q_��\ex�^�>7�ya��S�6�`]W��w8J�?��/�]�82��2a��F	J���e���g�+��p5v�� d�zQ�әt��h�%�ؾ]�ӈP(�hTcHYY�_�hjߊ����zTK3����VR.�������.�(�b2��J��s�$��(�?��4�܍߹k��c��b������D�j��� ���h�C1�4Ӑ��(u�p$�Q�ʫܕ�(��Qj[V�y�Qf�b���Q�j���)T��g��t�θ���lu�ԘS�ȋJ0>�*�/.Y�7��ۡ��P�IV��h�L�+/E��G=�~�6��7�T�dX�7�Ջ,�3�7S�E�dõ05x��� >��M�EgS޹2�hքx&��o�����3�΀w!��t^���"��b|��G�P]ی��!�I�ӱX�hѼ�����_oǀ�����:3�ş������_|�nL�cP4-1��x��t2#J��,�d`��sIu�O���Y����2â�-��T0U�`^Q�~������?��K$k��2m�{��a�N7***�����0����d�R�f[���K��8~��X��.Tմ�>?.����e9��@M��><0����(�a������>�?P�Դ�U����R�5)�8}ދP$�&�҄��sJ6�d�(�:'�;�Y"J�_��:0��s�BPD}\Mʛ��ٿ��s�S��B�������h]w;*�u��o�^�Ao��Nq9�1r��I�<8{��ܝD<�DU\}G?$'�/}�&W9��=7(k"%v�����	���,�a�-�9J]��o�5s��S�B|#Ô�+�n�¿Ӵ�Nxb3��i�N���X<m ��/���_�f�_��d���2�_SVz���jS>�7��x83
�i8�er��X�#��I�Y9���4>@�/��0eՏ�,�h��\�_w�6��K���G�����sd����Y���T�[݁���3*O�xLZ)�ц������w�@\��i왨[����ʴ���B	��(5*�9Yۅ�����e�,t
9	��4�9)98��%��d����-x��i7FR�c���|{0ZQ�O�%��y^�d�Z��YA �U�m��o2%�H8Eg���=��Wˋ���-jA�F&٠��dm�|ҫ��Z+�rt��&��{�*%��)�t�?�s3j��sT�����R\q��.%Jq�P��;�2�GQdY+Sf,�1+�������VL��$�v����o߉py���rL�i�J����������[�8��r��|d�|�����&�n[638RjE|F����~�,���\/���%��>����)�rb!N&�^h����>Ҹa���>�jʚ�E��u�ߜ�~w3t�)6�s��
;��nI�&k�B+�[���s;�x��E�$G��\�tg�E�9�Xd�p�k�7�9�:sR�7c�xƦ���C9Y�<t�L��R��4�(TY�m�d�ErzlJnX����vqE�ߧM�¤��_
�CjcU��?��)�Z��F���9e8��I&����7"�Ί��O�4d���$�6%�ϔ����	�OŲ����+&q�ÏjG�� �Xg�6�$� OZ;�<V�0�̐��Ϣ���6��z�A˖�sX��\������|u�]��_��0'���qiZ��8��'��cq�"�L�T�����PT�}�����1�D-��XY�WN2N�jK���FG��r�:�co�/�k$<��MQ��ϸFqWMk�<��n1{#!�N����~|�ӆ��*rw[=�{�,.M������X��;�� �~�y�zK������oܲ����F����qyҏW����Y&��@����{v������僸��N��85�A��&"1��}�o�/���fū��3.{�V�����\3��V���h���^u��@5�4~��[��v�GQQ�CBJw�{������h�C��]� nq&��/���	���i��۾�D��79�暑)b~d�ZY��~�����=r'��{=~��ױ�wX�m�b8o��R~_�syXf�ya?��7I�W���1���{qcg~���xJ�<�$*����AyΕ�-��/Wҗn؈�/���=nSף�Ģ���ٖ3��W׿��Yy�!���,E�����:�АQ�����f�28��V�d�[8��p�)J��y��$ �ު��CD"��f�Z�vW���Vly
���Z%F1�XC1u��v�W8�~����~���Ͻ�?�м�U�A��P^b������$s	�e���G���W�ƍj�S�Xc�I�RE�l����-Aյ�9vQ�X_
+q�xۋg����Ŕ 6f���5�5�J��+��ɘOo_��)�w�����0Z�|%%�������(--�PJ{�lۋ��!�1$g\�4�*�E1f���uO���Ҳ*T��(3*���+��y�6T)낡���hQ~2O��H�s�"���f5��ֹ%>ƙ��ۋ_�Y+����n���*�'<���5�2591(.�&X�����~�
����qD����FYi7�5���ʛ���j����|�<K���	��*�98Ԕ/U�iH�&�Zy4�L��V�(#*'�[��i&��Ab��E��ň�AQ'��VM����h0*L�\׽f*�?���N1��Мd_��D�~����R>��5�Z-����~"q�,�����*��G�Y��W	�=ј�r��o\]ĕ�����#%�ۧ�j����\������Nq�;�+�k�^;x!��<b� ���w��FD�w���j��!�SJ!�S��&���p�\r��b�0r�8��F���p �̿P�Œ�}]��'�L�;�O�O^: E��2���s*��s��)3����3�"��R���aa�o=��X2�� !#�X陚r;B�c��ӭUZg��/J���~�������ij6]ۂK!~Ef߽�M�	���iF����i=ʕ�ŕ����F�O�r�!<(����F���Sr��Oѽ�>�W��g�TO�����x5� "��`�(k�ܸkj\��{��o�(�$z��#�����"���	qEP��z���^%�cx�L!�c�siǘ�SǑ���Z3��Fÿ�c��C��߾ye����ڎ�^�>�<:�߆R��2��q��k8?>�wc������?c��<���H�qT�[`4[�c�7��kq:^��!j�ݥV{?���I�|�
�y�mE���H��6J���P_%��R�E��ӣ^�I��uI����iҲ)��7u4���J�E��9�X��Z�TsL�����E�N�@V%�I��}�d���^�Ӝ=��(.����Yh?O�=��d	�z�[��'�%�8�<���6Yzz�KKG�2�ej%����Ĳ�P���A�S'���ރ?{�Z}�/n݊�z��]��XU���l�§w����]|lC��q>ea���rO_T&/E�s�{���|nZm\!��1X|'�Do��BAԍ���K9]�ɚfĸf8	���(oG�xnM�C�dM>R|G��4?���Qu#&���o]�v�Pщc ��{{ڕ?��ev�I�$Q��k�'��`��W^;$���߾s��MW��c��i7���tʹ�J-5;�8�k��eD%�0A�8��R p����o��]��z���ӆ���W�ʭĘ[�K'�֮&1>�R��M�P��s�����Y�WOH9�sA7z*�7�7����S����,~A9t�Q"�̸A���UI��Jaڔ����٩^|�|/+����m�老C�4��k���"�K6�:��p�iW��\�N�0���C9��h4gR��aNTR�OVc𬴰H\z���Qlo�뉦0���p���X\|!��_}�Q1|S1�޴	�����ӧ��W�Пb��B���t�)����z��t�*��2٣9��8Y<h�=�[4ZSb���F���/����h`�ɋg�Dw��Dx�| ������и��ƊM2�0]���0=� ������_�}5E''��G��C$�������防×��rv�����CI���58�(�_��w��>�DG�&Եl��dE�;���c2�L4%�󚼤���^F8��)�z� ���&��"����B�]��7���C�B��T��E5{��
e�"U�_�|�I��k�Veб�V��:����]Ės��Do��f��dF�-�O�&�u����=���XQ�Z�6m���'0��⥐V�M��*&�8X�z-g!e1����eI�?�m�]��[׈N�2])}Zd��cJ�3,O���k59�3�&#����5����7���/���^aƎۿ���v�DZ�������a0e�ج{����^�6u�m͍�E�H$��Q�����tm�7���ވ1�@��fl�D,��w��J�+���l��z�2��wN������)�͕I��*�m����������X[�߭�"�=(1FCQԖ;��c���þs�U�C��P�����TJ����醵X۽M��4.'����R�4Xp�vZ��bkV0:epV���nB�)���8hgl^)���Pj���ޡ���,:���[E$/r��Y��>���������Z����YPJ������|��볜��o�$� ��{q��p[������ee9Y%��c�*��
K�%�󘲜��l�PԠ�ݥ%�፼��UWUʿ��*yA1�Wv�Fc�	Ix�p�����7��VL������(���>"����S�L\񅋹�tZ3|�[��Y/��˹�C�tG�vx�.�}������`�
&F.a2�G0kE��{]+�V���a�����lZL��3n�\8�r�ҙ�bJ��Ă��،o+S���ݿN5Y�"a�N:$�&2�7ٰ
���}cH�,�eL:���u"����զ@C�n�	fd�Ǫ�{�N��������^�V�����*�W���ɬ��Š��Mba\�R�3�N�����7 !��:�^R������bV��ad�^J�+�`m�m�P/W>��6x��Mh�ڦĔ�M�Us��>�]T�i�Y�`*����ѳo!���~�t�����C����*1.-ګ�9�yCb����c8�����ء�'���)�c8E�3LQ��h����<?���=�L3;y��V�0�!�vI�O���L\Fe��0蹂��^<�U�����qb"cŭ�Q4�	��i3�\�9��.^�=e9+Mh�9�"�!�U�j�����տ7����\��l�t��X8��0j͞�ՋY�+rU}�.k8e���f)/]4���E��O(��:�� 8;g(WC�_ж���c��C'�F*q(Z�cN�x,7U�=}�	��?`�]�ȟ]��YJ����\�!�+��=��4��X��w���R�%#܎Y%�T���EKQhCX���O��i��.��u�Y�x_ؽAV
����B\����C/��T� 4O���h�Ӝ�N{ m��0�E���.�J�ˌ�	�3��+qE9B�T68�㯝x_��}��-����Eh���G�Lɂ�^�<�BWU%j6�d�"�����i�����n�p�Gz�j��� ��w0��8ӥ�E��sm�m�bE�g�g���I_�KKB1UeNĶ���a�'�W�Њ�Ez��v��+n�U����ӽ�pWJuű�	iN1���1Nhf
!�E� <ӏ�ou,^��� !�i6�5o��H(?�v�B{�^:t5�(�*϶��|[�!y�#b��Sk[i��'�i��б�&ɏPtf3�9�&L���_��I�ŗ0�:c�Ç��jl����؈HD�bd�Yk�n���=�3�r����Şz�rGs��CҴ�8o��������-�MR���֊���d�bc���6�uXR�"���K2��'r��,b����]�ޟ�K%�Y8A��o�;��3�;)3�=���n߈Dx������`$�eh�؂�u7�F�P���T�;D���OC���K��˥�A]�͂��0���Ӳ�J$a�|�� O��f�U �6d
���2��ě������]�]���|�Y�׭�4��C�&�mz��rg�nu�C�c��vIg������qɂ�r���Ȓ�<�9��]�B��`�=��$�&)l��BQϝȸ�VU!�bN%u��*ڱ���^ZC�K�B׮}��pZިt�1�n��5ɰ(�b�7o�,���К?Y*�r�\Y!�&�����7%��X��C�*"�-���C��ݒCg��rǽ��$�2@�bQ6�t�XGt(�}����,��)�3ׯG�R��!TF��RY��i�k�����_gBk@ �Ƽ�@��z�ח�"�P��� �A0�A$G�g�ZC8;�Q�����d� ����a�e0,�(T��7P%f�d�:�d�1rJひy9�2>�OO�j�35I�g�߫VL���@q�ʹ~I�2�lf�~8��׹E���\JWcؖA���6�D���S�b�(	�@]�"j�N[��;�o�,<��1<wb��E��AS�z��:�^\؋S�2��b��h���	�̿|�&��Tc���A,=����<j��H�ܪV_D�����B������!E�>��-x��9��bI�r*\8(J�r��i��+�qbԏP2+zc4�P�c ���}�e2�u�RY�FI��Ա=�R��狪kJW�ҝ��'����cM�w�N'*�|E�׺n�,q:�"v
�ѡ��?��_�T>DDq�D�o�����G��D�	'1|i/����R�Uۘ{��K�����s���B2�ŗ����L��F�P��TΣ?��Иbʬ��Z��U|�y�i1��������q��f\�g� r�R<�Y����JN[�6wwng�Ą��6��O���0)E<*�n��j���ܜGu��S.�JY[g�#MF\
��S)Ԋ���\��J��E���F�m �O���&8�͢�~_ޏ�}V�T��̎���������������P�I����9��:��QD�c-��ڍW/��̌��X�L�V����9��^���������+-xl��D���lbQ�~eĀs>,9(2���wYQ���t��:[���98G��ޅ̒"P:�յ?�aC�#���
��/�)�}<~�$Ք|�=\TFC���PրoxZ���6�_R��"��������U0L��1DS*�*�u�ƜU�/ˬ�� E1e����<���mk��)e���ӂ�λ�51�t;��J�e��Q^�Mq#?��u{O��u�c� U�3rGYu�Dte�u0Y�72��k��g�6�-��$�D<P ���"cJ��`��'˟XֹX��l��
u|�7u��b<`K5��`�&q^&�w�����)	�Lfl˴`[��.�hΈp�
�h���e$��iv�a͔�e�:򕔽��Q��2��t!�b��,e(svA_�LR�$K+��4�b�����QKiC��4��D-���q,w�Vu�f{]����)�({�r��G�asNnOF����=c^|9�|���hɂ�=��dMI�bFYok������~{���옪6^���W8N�l-W>;�|+�K��2exH���C�,�Ȝ�!:��>�L�O�3�ɔN(g�F!+��2HEF\���=W��
�������sq��e-q�7�[�#��ҥV�n�u��h��ԗ9LdK����倧L��1��a����2�D�dRQ�Ux���t��b�m�W��fK�&��1�8��)�E��L��R���3B�E��{�v�b[y��*e�*���rh�c����×�������M�T��hi�(u�Eɮ`m ����OH+v�]��!��Sk:�W+�L�R�{bnN&�G  ��҂�]h/t�f7��U�Õ#�4�嬕���&p�o���+G�1�)~�=���ʱ~���j�fC,��ӯ�y���p19ϦO���B��AX�a�n�)+�
3FKQ/,=��Qq��j!�Eq��:�^T�%�G6��UE���u��s��z,�z�#�q�7[��ժl�ڀu���>>c,�C����P��7�m��h����Ƕ*#���"FUZ�r��vJ)�{���U�Ol��~�X�)��9g�G2���R=��(��zh<�����V�U���uk�N���X|����Z������-[$V��&[����#�+Gwc6����_ ������ �&���x+Z5�-Z�6��в�5��������Z���k�.Jӛ2a$��ݛ���=p�l5���Q��%��KP�&���~�f1�mW���rJG~e��a����yv{#�\-��b�k��g����=un��͛��ы���S����]Ꙕ?���+����]����8�*�*�p��eƬR�.�o4[��=��I�,�b�Ty�~�����ֶ
��3�/�Đ[:�
�ۦ�ei��C�DH�'g�X,���aͦ0�G��Z��5c"
�3�����	\cv���h���h(l�\q�E'��4��R��$:��+%reT��b�7[$�+�My��P]Qt���!_�k�����ա5�O�:�p�[�L�/!��FB@�<3�7I��:5��q<���@L���K)��I1Eo�  ��ҙ����V����Dc�g�W=�U1٬<�d������5�2�l_.����b�I���L֢a`T�q&��9�,$��Br.��d�h�ٞ1���J�psG�o�;�?�����$j:� �S/�hV�'gf�&+�c�,��ݨp*g�l���
I)�=t� �$�ZC��QȦJF7�z�VJ>EY�J�&�N{��u�64��m��14(shp�t�@ ��b���i�6�J'�U�	�T��H<������Ԭ�xl�RXJ�i	��:W?���粪s�&�^���\�S�	ß��n��/U���èm�H/1�9̬W�{H�l�\x C�R��Q�B(9�,:6���)E��B述��.��pK�Q�����XSf��_V�.���L0�+O�f�&�#��Y/ȝ-��$6��)e�D� �a��� Y��[ެ��\,��!���RDLd���x��blԤ������;�+�d;Z���O0�Ƌ�Zt��`>���N���+��{�w�U��*ڷ�,r��W��=�mV�� �.�J�Mf%�|�%���i�(X�u33��B1B4� �/�h�w���d��WYd���Bf��b���#{����DFrKβ�������I"K`�����\ȿ{�0o�6?If�t��z�g�S���JY\�����<�@���ʷr�"E�86�i��~Ά.�������Vt�chS�#��2帐l`��:+�Ӊ��q�I��`x�d�^�թ�,3���o�>aN�Ъ1E�p*�౦�u���hn^�$�q���x�~,���C���G���$HC3+��8w�/SXg���}1���66�*���8L�D�������7��6���5űYD�s�l�Q0����.'����b˼"Kj�a�K/��H��ł�CO�c�ֺ���H���z��ڗ����T���͢T��V���4�
����^�+l��0��"�0�8�79�(wYar�Z���A� W������_�,ZƐf.��c��7�U(�����3��CgD�)�I�z�V�����rnqxQ[����us<V�L�Z�v2M��2«���˩q�qD����$����^��a��t$��LY�W1���a��J�h4��#�)����<�i1�!�>ZE���Q��#=�!�:ϼ��~�J���&��X�IӮ�¡�Щ%�� lo���8�tH9>�c���R�C߆�FҀ�L�pp�_���:��<
gU�����>�9�*����`C1�S��n���g[�|�-�}�e�q�b��o�?5�g��M���[1|r[w��|.�1f'�MY-O䃛S-Ҽ�Ǉu��y�b�G����H��^<X9��5%�q�?AYy�Е��c�]H��\L�q*^>U(Ǳ��GS�:�7�G8,F%YL�ߎw`�ĳx9\�Hƨ����۔�4]��KoD$kn>Ih����[�(�0K	e�_���]j-u:މ�/;���ŭ�V��H�=��b��$Ƶ.��a�=��5�	3_H�n���ـ���1yH�QR�2�P�- ���L�(����i�W��i3�A�P"��@���!�o^\���<�Z]����%���XY��"�2����R[�%�+`�N����1I�V�)��!�҈7ϭ�~p�@1UX�rg�������)�e�]���d�3�5(��8���L�_&VڌT߳���-ܚ�Rf<�(��Z5�E[$XW���h#	����b���4�Mݹq� α��Wvo���������J�Vo�}�a��"����:)�(��+� Բ��<��XDb�RR�غ?����y��������E�X�1��(�yA����`DĐ3�����D=�Fu���rH�ɮ�)�cO{�0����J#����C����+�,W���4T��Y�a��a�a"m�h�I�7i�����MI������S�K��Bk�#����c/�{�G�|Ӏ�ә4z/���Cx=R�X� ����n!pu�]�����3��J�'6
1)�v�℀{Ԭdn��'/���LtwL�*\m���{g�b�0Q,�  N\��7#5�P���йn�˵�	�w.�}�G��n�m.��D�*�n�A-���՝�v�F16ч��������F��P�ݻ'����ː�,���g��	e�P�g��Ր���@�.�UIk�+���UD��9���x�j[o�}��,�m�,�-]MJ�W�J9���>v�m'.)�A=�G�7�~��U4'���8w��;pCď��c�26�5�Bܮ�. �
 ����h�RC���aT߮�j'/EлWF�|�_�-�.�99�(��Wߠ��.1�	~��Z�:��URB�3@��	I���Jq �!���Bk@�g�Z�p�Y�b/̴�)��_��z�J���	��Ё+���͝~�]��J��±�N![��������CP-��s�]/ K��5��e@k̎YM/ւ�W���?�KϜb�}xLT����|�g�nEC���+���#�D�u��N]�Y�1�k��J|Ɠ�$p=��ްH��ݎ��_� q��4���kd�ټ[��߸��
x�bA��1��*�⌭+��! ����g�/�ļ���Bt���dawV2J���+�|����֞��r�U��Gʡ2,�8���#���Z�
�&���tKH�
!O���G�|׋�Nl��}x�ET<�͖�ͥ�X�"�t����f��觑Җ�6� ��պ�!ZY{eǴE�+�~�su�EY���Ν�������_2�q�0��ы�������-�8�S6�Vc e�_��78��u^{S;j�7H���3�}'�/�ꊡb]!2/N���\���>L8U�?y�]T)�7n�"���hFGk���xꩧ099Y�+++�����+�����׊"
���)��a��vE�ֹ�u]Ҳ���]����V��1��Q>���u��X��n��O���k�[7����0��㭈[������Q�a
���~�$�[)�a@�+�a�QS�S�\�R%3Μ9�o|��j������OJ�;�(����$�3�?�Ww��~z����Q�ǽ����(��i�i۶�]ߍ��a,m�p�D۾�'$Oo*������w�\��_������k8s"���O\�������7!7�J������7��p�����<��s���i��� )�ߵkWaW�k_'�A�yOO��_L�Bi��݂��� ⿵�4(f0��O�oS�6�_�^|?դ��z��:���V�ph���^��Z�R�o�iJc"o�^p��޶F`5�E���W�����آ�����?ceLd���������Y�W�փ|���H��z��>�\p�3���P�V#�8:�2�5JK�P�&{����@������g�ޥ�_��}�ӛ6J(��U����B�����Z���L�0�k_�ȼ�T(
_����c����
�4��b��@���MwJ��<+���Z�;4�.��_Af�-2�,�8g�`��}��0k�)�x��#<��GrR��DN�ʏ̤�cu-4�VV�Gd�eMUUUappp�UB��쿦��X��i	V+r����2�|!B��`E m���E�7��ꢕ��{�Tߍ��3�58��ح��{� ���V&������� .���G�l�b4dQ�,+�I؋���s�ќIg�}���Ʊ�v]�O_酻�_����eE�=���۽�J����!8iA����k���'j\k�Q�W����GM"-�˕�w�(��`��x�b���D)��a:�"�1%���hҢ��}��o2�����ۜ�̈́��v��!�1���AF�� |3{���K��|�wbxx?��ϋ�.z�M7݄G}t��^N��9/4a�i��J
���p���#��?���������(�ńcn��&�K�j	�=��+�D��S����T�n:��00&�d���XNށ&_uY��{�l�J��:�b=.��t���/~�6m¾}��U"&-+2Dg�jM�CYc@ 6=���6�/�Î�1���NEc)�r!jq�}�9��T��	wv���c�Z�g��2��fހ�5˝���lڞ�(fL�p�5߬��v�ک^����:Oz3�b��ly*�j���_���w%s��Ї���T��ճ������W@�7/��&q,}p1��\��p)O�"9C!�ϝi��hRΧ�݆b��Fl���G�-1#CY�|�����z�,c-d
V �����癎�.�j�Р3y`؋�}12\�GD��eq�(������~FciX�ׯ�[�����e�{���k�����<tn,��Pl~+IK�-�?�	����!��q���s��;s�Ϯ�Ϧ�!#�j-o/��h������X�$�x2��ϫ�N �\5�+�\�AQUmNcsIPk�)T�m.>�d�r�5�Ϲ��SiFUm�R�lLE��?��p��x0E	K,T�vK�e��P{��J�-&]w;Bx�r�5�p��H.�31��W���fAǘ������Ύ6l�� 셃�Y�x~�^EDY��lP'|hK���D��%��� �~�X�J�V�K�����c�l�|�7��E��>�����˰�8���lW֬IC����𣧺�ozTy�%���j{i�wo��X ��¥d�tԲ-����=tN���{�2�����۰I9�1	�j�KE��	���`ݖ{V��:l7_��~���1�v�:�rYc��e7JJ�H9ȁ����X�ؾm���'o���3e�"�VX���2a\����l�d���g��h���bM��m+��W���_�]U�ƶ-X��^�D��J��,�2�@��k{E&ZJ���FV汶�ag��������s$�m�H���9����r��S�3����)��S�^��}#J�����'t��� e~v[w��t3�����v�~q��m,�a�u���*�&7����G��a�6v�s�A�dLJ�gfO$��5r�#�Q[�1|��Q�ǐ��H4���p.n��.L�hF�6��k9��_�A��q�V��z�uf�'}��l��,Cs�!Tׯ��U��J���*Fч��	����K�İ*q ��г��܉��v�	E�>]|gGF�R�]�����u�q3�DH�_V��?<�ӣ��5���%m��^բ�����Ѳ�6T�DT�Cj���w��ρ�`������n��n�C1ČH<�s3~�kQ'���k���~ǉF{QE<s��:�1:JC�!�L[���6<��/�C8J�Z�0ǁH9�6	��HH�1�I�K�nͨd��()�<�
�K�5�����w������qZ��}2|//Eױ�_���ɒ�j�'#�:�,k�tw�bk�׫~ȼ��Ϩ�#�4B����y�P���K�tȒ�T	�S�n���Z�����c0��x�+�� =ߴ�:/CX}�'=��f�6������Q$n{y�ReW��d%C�+ѧ	c\j����]u�#�Cs
�?0�̸p��/��I�������)�Stڱ^�ڔ���Ѵ��iTd�Dz�w�It�J��,
E=8����I����x��P{$v��!�tf�^�g7���+�<u]��Gz���Ԇ�T������\.IIO�<x7h��z���aei�<s�Z�m�4�j;��F�h>�*j��⫞6x���£g����p�Qb4����uU�����d��L�E�:e��+�V���5�4~���[[�v�G�#C���Qye�\
���q�#�]l��pU��(9U�l��[>�\�	ܗ��?��e&0��ZV��3�ɖ�g�]T��2b�>�#S�zl�z��9X����8<8����詯V4|&���Q�nQ��$���)e���f�Eo)	�	���`V�s�ҎQɶu��g��4e�K�J�s;zP[Q��>���s��>c,�}\'����-є��V�c]]�c]I��w�b+���)"9�����B[�Nly�bHs�ؚXN��h1�����z��3�\n3�a� h,�
�MH���lҷ]�}p��}\�Pu�H����^p_���~TZ�(US�^���ze.�mya/��Ӝ �b��&nB)�Xt��F��2��c���}tk7+�d;;f����K��*!3�+fX&3���L���oՕ��ѮV����DJh�G4�GM�\ e�3V�
P�t��d9v�U��F��e��Ҕ3kfY�>|�(&ٳ��$jc�����L@�j��j���Ud
u(q$�5�
��9�8�؈C��5���^6qX�6�#A��W�/L��?ލ���ׇ�C?F���PQY�A�&b�=���O�P�@g�&��u��A�`�c����^���Ub
�zϟ�"M��[&�1\|�4^�Ԡsb �������y�^\9�*�Nx��g����X��e~=�F8�*]��(Mb����uXj�f'�^���;���6M�:�άNrj3�W�}�S$c��{G��g�zE�8�%�S8w�I_#>�;���O��Z�!��8.3���Eh?/��Hʆ��l��H��k9�9��DʬĒfMh���ݝ��
|�f\�k�St e p�]�RH�P�B6�B����ԗ���x��uY�F��+�`�W�\$�Ơ/�~oH۳o���"3������c���r���n��}U6���T���Pq�u���63�1�)�YՀ$��r�/R��n����F���
b
��}����3E�w����=���=������Ug��f�>V�)z;�}�]�����	q�Ãz[F�;����AUU��`�WOS^��~1C��ߢ���˽�a��mӰcF����������W��']>tt�@]�1{��!��ߋ�	F%����2�D�Q4&,���}����9�~�Lѻ 8	�=��s��{{���p/ܵ�b1z�.c�w�����jf��\NkKb��Ӌ�7<������ΟT�v��qo|C)��"������	�	7�g-����1�f�C�2�"�0��F�6u���Wr��Q�}����U� v��%�����^"\WV�"����$.U޺cf[�n��Mݲ�[$F�P���I��]��.�O�]%����G�/���V�b-ҊbY4f�c�L�m��Ռ���H��ַc�소���5w*4�r*��c��]Uׁ�5۰�wR�Q���Z�pմ���� =��
���*�	�%&T(���dW�)z�_{�����}��)�'|2I��[G�[w�D(�h�EHj5P�:����*��jE���\ e�����f: �t����V�d��W�u�&��ʠ���k�kYJ���},�)��?:~Q�x�R��p�O�Q�J�^H�-
ӛ����Ci;<��о�X,VI�phP���D"_����Vua2���X';~)��3���P�<��K� Lgr��r^�o��
oڌ����o�)�Ks������3R�5H�ݨ�'�Q~�5to�55�i�-�}g0pi�lJ�D�ָC��mM�:ᙖ�I��1CK0��A|า:��GtZZ���Xچ��8ۀ��(uh{{��I\<���{�?�2H�\z�߀ϞQ�\u�h�����˾R�:5hu1��YlM	G�Ɋ�E�Kuf0ӧ?Ňi,��,"S0�H�J��U�d_ĉ:s
�S/"0q	�V�;a�wx|O������^~p0Z!%�7G�hzC+&�b�z�"u�,b�u��Ŋ���|����)�=��� WY}M=��}QN+1Nѭ���l�N���A�@��|T�DZ10�3B'��Ja<k���-�Jʋ-+;h4i9�w���ae�>���y4z��s�11���t�A���e�(����U�<������Y}y��Kv����`�C��FUV��"ӽ}E�}B��E�ď�fdS�w�s3�j攼�c���!leЙ���7�!��U�f)��a�^h=��lX҆Zx(&d�7���|(��3c�b��+�G� P=�ݸ���  n(�������;�[��MӢ�������Tb�r��ʔ����J���0J�9!���!�'c]Zc�=�ϻ��U[����ط"�Ğ��x���K�ja���#���mqUH�;�}ؘ�Bf��/�z��dZ�~��\�נ��S����=��z�׀����l��W3�m؉��?���Bo�:����2Y��Oy�̷��mkĢ f"+�2`�ޒ����)+eFn����D���{�Cx��Ö���kg��l�����x�e��x����h�ޣ�Tg}�0�"(Ґؒ�Ծ��8n��	e���oym�l�@~����bʏ>xLY!3���o�*@��xR@A�����	���s�b�.�b�"d-J��ݬ$� n
��3��۔Ψi��٦�s�hn`U۴���i&��O=��-u�R�I�Bk���W����R>@L)2�^Ō���3�K[�X���D�͊ku�j�z���[��^Bܖ��ʎ��.�RLE�eD�ԇ5ϓ��+�u�w�m�h/�_V1�����1�*���a�\H&���{�}�M�s���܃�z��J��^�@;7W�FÅ���
x���$3�
@ʝM��7��wL���P���D{g�
S��L�r��KW;�����n� �$�g�
j�Mu|a�2ū��-s��+l����'�ҾY��ӆ>߄ )��g5 e�o�Z�"�X[�����T�o��f至��̠� �:�J�d�Ʉ-W�UӅچvT:5h�|΀��s�?����⹊�����j��c?C$8! �&�YjPG.��#�a�nՊ��=}E�M�sc>�2�=�	�_Ly����s���E�|����qSG��rz�'�B�u��߇�c��ҹ2�>�\9��}v�N�ϭ����@�rT��5�����$�S/Ë�VD������.��o�=�]o�\f胢�m	��5ؼd5͌�����&�5�&*�F�N'���Q7�F\�#9�J�Ͱ��N٬�����������h�J��bJ^K\_f��Qס�F��Y4g���xY�n����Wy�y
g�N��^\  ���Xm����y혱����9�T,��~E@��;H�j1�:3c���� �l^�y�㑿>u��k͔9̸~(z}�NI��`) e������4�Ld삊Q
}��Ҷ�˯.Nֵb���2�̔�[u�x!��@�z͆,�Q��]�?����4�\u�[t(�Ao`�q.>��A�V�����c��^�r��KpS���|c� 3z�Q<\9�.W)\�	�x��8����&�xF�!�d�<��oh�Ɔ]�D��^�v��ϼ��3���Vi�b�Hn�F��C�־�Ɠ<�\'fX��y��fIK\�q|x�m�%��Al\�k�܋{��;����Qz�"��i+��Y,���̇�UVl��s��V�5��;>�t2�{��V��ɔPC'��!+��w�I�*x��u�������$�:���R��n Ʋ����a�[>���l�����'���R���F4�-���z�zz[4�c��u;en�Bْ��E���5h�]����1����+����7K���d�O�� �!S�
+e1�\g�a�}Qr�X��ڥT WHc�N-��� Rv���ܱ�_�[�*�ܬ�|�p�j9U����p��  ���[L��R9>4�-M��%����u��]�)י���\���A�I�@k�)��IH;�z:�k�^�0�(��A�E0�Pp�h�d��Q����2��M��>�c��pT�Ο��#� �|\7p̅��~XSm�_4!�V^���!�0!��#�@MC�\�(�#�5
�r��k�L�R�5&'v��T_�o�a�D"���p)nC Ch�,܎������H���1�ܯ���=5[��i+@ʷL)S����4m	�\ӸN�[S�Q���p�1�G�<(�@S�`̉��l�A��{�j*����/��P��l��|Ѹ��L��2|F;��^�)j�����-�]w?������!��kCO��|(Ë�Zt��`�����,?%���g_�O�b�s��Y����Y9���~�r����h �C<�Wr���j�ӓ�K��c ��x߰|ɔ�ĝ�ȗ;�;�"i�-�C�ۗ����4$�Pʆoy[�k��]8�"�B���mx6�,�7���$�e��e���≩�0�q�7�@,k@sIF�����D?��쉬p�o��7:#��a�ro��h�ڬZ�e)}1�n�BkmK�����<��^:�l`U�'�e0?@"����4�>�yL�D9�L�^�D�5�?Ĝ_Ӿ�_�1U���h/����A_�Zl�'g�Oۛ���lnVG3�]=�i5FV�$��U������w�h�9����^=|C�q�)+���ņ�-�,�d
��\ح��.�zx��\�T~v�Y�1@���Jv�R~�Ý{�񦲹U	����aS��ɀ�Ю���_�Y��ϸ��2Y����������4|B��.SJ�Ɍ���5o�PJ���
�8|������R<+��@�,��̠i�Ж5bY�y��Y���c
I#����o�gv�`\9��D��"h6��c�ϟ�'G<�_r���7H�ڲR<����?E�]e)��=�����¿��ݲ��~�Ox����n�G���l>K��cI���	�yT��Ns�W�csi.G�L�qe8�v�Hu�wCx�5�{�S��t�rd���!�:i?����uO�Xb���o���������.�޽Hp1���R�Yf�"K-f1_8{��_�=i8p�r�t�a�����A�L��g�T^r3���}�������g�c��~z�����=x����qebS�2y���t	���s;�_��Ƕ7�n}��&���;��c/�=4"!x]�C�Й۝1l��WP���e(B��^��JW^��MN���F9�;�<�k��.�8tfI�K����V����}xt�Z����⿾�_v��$�'���Aʵ��:��C��b��f�6�Lf�y�"�y�W��uRA��}�y�w�n� ��}�L.yø�9�͵e�q�a�W�5�7����W��A�WNE{9	����Բ5��;J*e!��	�۱�vl�>^g5�ey3LPj��1����YN4��M]�Pb�[����[wsG�݊\!,I��O���Z�+�O�{{�%w�
C��t4�5�O��m�2�o��"���:��^EO�N\���cS�;�3���XB뚏�TMl��+a(��:�5��މ���q<�!����-�p5ʇ����YlMX�,W��e?�@�(������K�{��7�yÄ�����E\ڄ('����ch@Z���b3��x!mWh�� �x<���ާ��-������T�g�WW�Gz�0����_Zp�P1�	J1L����58uɇr%��uT$]u�0V��a���ڒ'R�T*,�I�Y�=���˙�LƑfy��2)nnh����]yp��y��V��iI�۲%���q0`;�i!G���t�L��@�N;�%%L�@��@���f:@&!)�6q�����6�2�й��]+�n����Z����dO�̼��c�����}��}^�H�t��}�,Pm$o~E��%�����*���7�:��^������"H}�]�{��Ú-�<�3�㟞8�}�5���3"��x}��.���n!ru�-��?�S��M�zev�M/�a��k�%j�]8ٺї����Z�i��NV*���Bw�����,�~�v�,�O�[�C����rh�a�������B�V���(�-�<f�&���/�w1BbS[U���a%n}g�(@��e���4ʗ�ӠE ���\��|���B���^v�6"���Q�����+�}>\�{M'ph��~��+�\*��y���[�������b�EJ1�:����,�,ǉ+�
���^β3�Ch��&��ơʾ��*@�r�#r��>8�k�Z�99y�ۑ�a4|�&���B��3C�N�b�9�bܭ8Ϡ[4�j�:�v��݆���p�_�5ř�rn*����ht��f�+6W�bIp]�>�,������g�:<&06A� �ٽ�v�#J�����ӱ���wM�8�Q�U"��xZ��y7�=�l��5܅~{&��\�\�W���#8�Q���B5zcg�ZW�s�z�_��{:���:ԋ6�����;��{���7���w �r�+X��/�`�E�PN0�߆Q�Y��WcLQ�^��Jۧ�Vb�� Vt�W#�s"'G��8�����]����F�����VWh}��m���aDb$#H h\$���AW���i�Є=jq���)�z9zO&k}F��L��v��|ۤ�Π�#�$8ۤ��	vr3�6�)8+g���L�Sv�o�r�U�2��͡B\�R��u�[��}981�R�턅�iο1\,+oeD�"�D��j"<��ن�r�<9.Z�U�HR󍩬�T�9�G8q4��f�>4�S$��b�G�wR���:�o�9��n���q�L4�����H搴�F���H��#GT7�}V �@���k�d
�����Ao�\zT��TK��u�E������T���M��x�����M�[�'UO���Z)��#�S���s~�(�4�>�ͮ�l\6��.�i8�ܨF�9&��=��Ry!5Ւ�Z�=%=^� �)����י�"\���o���<:Yg�>�s���W{���*�2��8�Ӫ2�h?���oFIf���Z��}���`��E��qP5���A,Ms@�a��{0*�(O����E_?nط;�l���-�e��&����kIi�=���"�o�B�G���xщCf�r@���R�0��FM����AeƘ�8��;>����p��k�sE.�D'#
;�{/�\�I�f�%�ıX`wd਌�sԡ&d?�Q(Hs�\��ъlȹ2�jeВ6~��=K�C�}�Eؾs'��b+���L�R���̬l�9�Q,�� ��L�/*4��
��.�2kw� vd��(ï���q�x���x�ָ*w �����kP�|c��F3�\<�U�#�i��\�1nپ6윫))��E�Ox�v���!-��x�	��L�b�֭ؾ}���s ����&��1�q��������yΌ�ЫLی��P5��B7��F��f�ʬ!��Ƕ��nkYی���Q|��[�]����Z�Ҫ�B�M�~�>1�����|����-M������S�`�`�ħ��f�o�EŒ���]�|2z����>��]}ʖֆ���t5o���՚}Y�Kk|����k�j1�G�N0�WqVo��_�1o!|"4��Ng
Y�I�/�.����l$�b4��EK�'�#��k�u�:s��.mt.�Z[S�]�b�,�^Zc�cT��n�YZ�k�]��D��u��/�J]��)��ʠL]'�6'g���f�/-<#��k�n�P��-h��ҌI�2����1� 7�5���ԍ�Y��yvfi5C	 3�6��KFF7��[V�d�²g��Tx��E �eɣa��'1���/n��ӷ݈o���ۚ�:e�-�sm�ǓV�5���Bog�R&�2���NR��v7�w̯ˤ�b���sZ�@�9��U�A�� �%!�3�m���|��'�H�Bn�DB�Dӻ��5P�(3����6��5�*���׭�ҍ��p��24v��V/2c��Ԭ* ^�w�\�ϾHo/z��5:��_wT��n��WX���v�7���Q��z{�ƾg���1��=q�=��Cݓ�B��r��p%� CCC8r��H_h���뮻�m䄑d �� ��7(#���L��*���m�H�� 5B�$�
^��O�ѵ�WlVe����4�?�����IT���������w�Wym����'�۞4+AYn����~]���z����Z���mx������ۃ�JY!{r��46����e��|�ǲ����-����5!#X�k6W���{��U{Y�������D��!x�%t]D~Q��Ɓ���������ٱ��oʏ;'3p���M��K�;aӍs�����ܰ�
?<|R�X�0˩��(��%PQi4Ӊ�0QD�����0�XH0�y�����ڼFӔ ���s(�3j�KOl<׻����[W�Ye�n������fx{y���\݄�SqDL|_��o��sǽ�n�6��Ki�R����*锠�	뤪��>�X� ��6�+��fK�E 9.�z���;�ke�it[�_`��.Բ��i~=��HlRo���r��ru����=��[�7�0�m��|h8�`��H ������2��<I��^�����XV&�J �/�z�E��[�S؍g$a
3)a���H���'�/�s5��ʤ�� ^��!a�]���"��V��
T� �#�z���% ��Du��F�d�&qQW6�K�{�E�₨y:[��3�����B0�z�!�P��� �^FPÞq�k�c[�Pf�
)7�rpz�`Fɒi��j�n-lEma��V��æ�-]㥁2�X���R�}�zT��i���n8E5d�U���3����`6]c����|Q��������VC��G������.���d�>���gݍx��MbrLS{��}RKkl_�v܄�lk�h@L��~���j!3�"���t�_W����;���z����m��ΡT�N�[�@}bX����K�l��:�^��vj�O����!8N��tUn*�C�w`wv֔`��k�������r�U���3ޓ��h�Kg.���R����7C�k�a
It��縃A�	)�Iy�TS�d"Y3��ŀٟۅ+6�f�^���
!B�:��|=������W�{�9aK}�se�v�����`����%�NTTo���C�}=��A�DL����74-�0��Αe����֖�x�=SVV6g�6���������؍�(��`�s�U����>�A���YT,�6��_M�,MG��cˑ.1Y\�l�Ṕ[��O���ە =�Q��z��&պX�YB�ܱc����̍R����?����9�R��"��7��kBc�I�P��|��Չ̴����)�A-�^܁�63�W�HY�7�v2շheR&03�������q�2;�/�\��9s=�DH%�����i$>�cP 3eܖ�p;�V�V�L�-���nF�d�&�O���Jw=�ZΣ��YY��0��wF�����Hvh]\@�Y�s�F�.����R�Ő!LP�%qg��9m�����aY\7��e���E���安"�!ZVk��85Z���2���� ���E��d:���A�#8�хׇ��!хr�z�?�/�r���J�BP�D���k�T��L�����.J���qR���P	V:��v�'��݃��%mm�������[2��)�}�'{���:�d�م�fp���/��]��ﵩ������d�7j\�L� _�J
����Qcb��3�lj���9�<&ˊ�l��T�l2@A����̜��4Y�6`������I�YK�]Q���Ƣ<�ٿ�T��N��_�J��4���������a� t���/Kq�[�2.���;Y��#<���{�~�ӛ0>a�y��Td;�� +\DxAD�Ud���M�R0����ĉ*�w�ܩ�&2��=�v�
�6��� VMM���oM�y� >�����ǯ����:|���زe**� �566��߰aCX{��*ǁ}�9q�]�c���*��[dG$>~*�C��N8��e�S.�&�;�f�G򔘅�i��O:�ʋO�G����ÿ�g�j��OW���E��*�(
%�Ya���>��F�~�i��W��v���Q��3Ϡ��ZG/�O$S�]�jՌ٣�a�����E�����+���{�w�y�>����s����#�<&��3+K�9�
a�3ٰ�<|���^�||8�5�}?`Ǆ��,�>R/��5<������9b���3!(3ΰ�HDr�e��8Z��y��D��bB`Xg����oy-���<�\���^��Au���Α���$\�4����	`#�KKK��k��"	����=/��,�/.AX�Y]eX ��&��`TY�611!p�� $�\�9>9�;�Qc)�uC,D�F�w���E�ji_���ٳ��`�'#�˄	ΐO��g�<#�Ҙ�E�o����E�M��J�S`�8#�/�} �I\"0�^*�====J�� Fsf���ҫ�B���_2'#	B�ub�f&�Է<%�Fi7�G�2��U�q�'�v�?���%��A[HY��#J\��4f�S4L#�+�:ǐ�L�0������o�|�D�قU�`\g		���$��\	b�?��Y���c��O���Q>V�vg7e
q'�G�c��Ĉ��k��i���\\� Dp*�=409�LZ�%�f�7����ރ��@o4DD���y�������+i᧕�G�q�'�C�K΢&Z��O��!̖���AZ�-����px}�}#�]�h�z9�YI'��MZ*��\��1�O�����>ĭ�aB�FsI�U���7<����yi���j!M���u*��E6w���ۤ� �E�Q�e�|�9�V{�!����4Ї"��%p�����1���)0�4�=%��+H�Hgc<0�ԜU���(���Xn�q��v��r�$@�='���H~�+�lND"�'��#o�e~E�-���{�X���؈(q-cL�]��^��Ƅ|��n�M�6�3��X(��+���3����E?��W[[���v�]�vzDOڐШe<�Dc}���oN�(��c��N0� �`�s-,v5�Dx�v���<�܍�[Y�!�hd���y�*q�1G�ƍ��SO���qMΐhGd,0���&Hy?�����~;n������}��:��t�k�g�)-C��M��
��$+fG|~W�s�?�2�"](��D�K��"�"'A��TҀ�}�QC��^Þ={�nݺ0q�	�o)�r~$}��n���ٌ����a����@��ov>�i��'&�ym�jݸΖW_}5&["AȊ�ĸ�٢�]]]��r���+�����L�;v�y6+=��|����('7mX�����Hnmm����!rA�DC5�j,^knn��Ç5J/�n��__�L�M���xg@��|����/��X����=p� �x�pNs/y5��"�Sq��]���E ;�]�w�x��򗿜�pT#4=���g��-W��x����g?�H��U�b�_ ��y~~~~R�׬ĺ�k4Vnf �tP�Z�f��p�'J7����� ��rd߾}ػw�a$�wܡ�Rq����~���l�-�ܢ-:�$\���j�����&OG���O����p�f�\"���/3�J�Kau�e ����$�]�,�^���*�,2H��o]��.���)�xH�X>��]�f�*E�P16�X���C޿"    IEND�B`�PK   �C]Yu�E88� � /   images/41553842-fad5-42b6-aa21-339597c45c1a.png|�tM�.l���$333���$�c��b;fff�cƘ���3�w�o��wꮩ��)uw��F:
WV�B�ǇC���������6X迖��e�������?�����8`�-c!#C�7������[��W����C��+���
+�0����_����7ؿ���g�l�ankg���Pvv �3�2������W�/��a�6����6�q_�0��u��fcac�ce�c����q��q��ͧ���E�[�k�j+��:�1��9�̙<��%���W�3w5x��ڻ�y��G�_�33�?B\�
�i+(���\L,L,dB�  @��̂O(�o��3A2+WWG>ffwww&wv&gKfV^^^f6f66ƿ�.���&��.��"�O����������=��s���� ٿc�u�+����e�w������3+���;���a���Z[�_r���L�p����XZ��������qp�	0������_~6.�����_��'�l�O)�;8�
�o�%��?��7s�_���Y�Yx����Yx�XX�ɿ"���ߢ13q5�?XX���8��;��/����3�|ڪ�.�n��7�߃���V���p�O��4�]���������'��$Tr�6�[���c�w���g�3��*��b����;-����ϦG���>?e���Y�0q'n�OO���`�N�п�P�X��i��G�$V�S4�FR���u�<��+:�3���F��$�ie���m,xx��q�؇�6��n���r]>>�.�-��e�v%8�^�?N�n�m���B�,	#3�o=���l���"���p��I�����@E��},!��Z���:��},���U�m��Fr�f�;�`��d��W�v�&"��h/h G��gMƳ��/+a�I�0�� i2`
�Q�j-!L�����O�|Q�����5)���9����F��l��i��`B�6���E�{o��H,�,1|��-)\)����r|������4_X���g��;U��a���9�z5s��6�l��^�At�}�b��Ŵ�>E4t�V��k�=�%�����G'�����㜠#��o���t�����b��� 9S֓M6!�r^�R�3�����!����ᗲ_q�$�';x������/>�S�K���Gւ�Ꝓs"L��u�����Q��ō�̬W?g���ޗ�7Y�k����$���K�={�*|���r+qъ ���{ 3���!�<H�)DڛD�{��+o|f��ߍ�ލ˗\��a��|,6#븒d� ,˦Pw���K���371� ��\y��6���qHdA��|O�:�I�?�0�$��ޒ����p����.X�߂��8ܵ�Ҧ=��}o�e�V�\�#�����J�H�նQo�kʗc��~�X�q��U�>�
�Mb��%
��k0�t���R����~Lh�_X���1'!h�߲B>82`��Py'P
�A���W���rv����|}_���U�X`Oפ���+���6FƦNJ��")D]�G��/L�7G�^v3�������5#�o
݆,��O^�+.�J�O�WL�b�!��$��`.:B$!JT�QLѡ~���rd5:6	7R_".nX
��j�3<Dl�4���#�?�1QH*a�A?�GUXy0Ug��Uv�!�/�"�T��e���5��-.�U���͇�_8���I{9v{���"h�{	Gb,��4牉�8��fR�bA\\N��a��e9��NE	iZ��
Q�q�R�k���Ŭ��>~x�=�ǅ�g�h~������WѼ��j�\>�Ք�1Df����C7��~c��ץP2�%̈́����R��~T�m�]jp	�^�z��S�59�u`R4��N)�*E�$Pe�z���LD2�� ���tk��D�BE`K�5W�7���7(�MhU��<L�I+㹋�GK��x���&�-7P���2��_��eF���:����HZ�Ȓ��n�X 2:Se��$>s�Aq�8SyH���D���`���) �Y��)�����������)�5kH����z��=zI?�<=�v7�Z<x��1%U���GJqބ�R��� ���zQ�*�Y��G�/b����}tzx�=�]�(�-� �⥠��ن�2c��$�<O�P���؏�/���h�\Z��KC�\�PN>�;�&�/�nZZ���^��ׂ�HT��YJ����%7sԟ�>|W���d�a]��*�^��d�VO��嚬Q@���e	jb[gdn'��7����Q�\�@Q#[��8��^̝h�4q�5���8iXP��B�I-�� �2�⁥&oTАdX���0}jj_j9�~W�2Zi��� ;��2*;cjU�p9\Ě2Y^��`l�uL ����l3T.�ꨳ������G+,A�mͶ&?��&���20�8� ��tH?��1���%�" ���%#��=��j�v�W� �\s�x�H�Z�*��e��=c���_�p0d�i�=��t��I߆�
j���	A����b?���X�/�UΌ��]�v\מ� �+L��#������8o�򱏛P��>`�����m��,@ɑ����f��V��'����]�K��m�l�ۇ�����Q��6(����OY�'�7�SX�E�.��1OE@�$+7TbEI#���9��QjlG6(�����#��E�#;��-����$ƒ\է&��L ��MA7p�45#&�ت���D��!o�k���wf���0BKh=*���l$e�Xs_���\��#�ثg
� �x�q����VD�������C!�c3���@�p��Q�t
��"Ċ�Ƹ��ղ�D8q������z�o�?l���#tK�b6�'���E�ٞ�?�p$����6�`Q���a���iv�����-�(g�8��"���FP-1z��[�(t/W�[x��� g�� ���t�}e �|e�<QP�0F�ތ|����.`h��ln�����vEa/W�^��&	,��P��x�^���#Ӣ#e�/�x=������u��'���c���O��^���f�"EG�Wa/�R�b���&���@�@��W �~)��"JP�ݔ~�X��y;!n���"b�o����
�W�>_8�7_���6!�|���s�0��8=�QW� �m|�u�{�5�_#��z.- H�c�9t֟#Q�$�Lڟ��<��ݮo8�oUs[b�m��b���ϊk�e�˰ܑRYȐB�iI��I�"����&z����I�\\(ľ��|<�J��w;jV�d�9v<A4:*<V}���.Қ��sqD8XZ�
�����^`X�L1kC|��G���%q)��.���z��ϳ6X���x�8��/:6����Ѣ�lO�T��)vuV�|"���u*�Y\I;_˕����W��X0��	��ɐwi��,!��0���Dd���è�L�Sd���j־�E]��Hr!�TNҾYq�:���*�@�|���]'�Ӣ����n�?f�T���.yʭ|�m�~�Fg���:K=�ڬ΀��j��\04�LI�=:�{5+�~`nb��?#.�_����fd^�֪Y�V����-�O9'4���>lZ`�@��\��dH�9̚%�kPR䕢WS���P�RNe���3{� �h7fV�DkI[���U� v�2�~a��!��e����ӧ���qCzn$|)Bn�(�S������7�W�(��]V�rb�)� J�N�gx���T}6 �8v1��K<��a�_�$ĨST��!�ASC�%��3�S3�Pd��~r�'y(���$8a��w�o��0�t|�d��ҩM��a���Y9�X%⏧�W�����S�\84#�p��j�	�H���t0?��❣*���$G�d�f���;#5g�sb-�ńÀ�+ȅ���9�Ky���t�⁥�N�� k�[R���傾,jma������ZT��q"��<�9t~Jə��oւ�dZ�����!02�uÁӛ4�f�d#V���x3�D�bˀw��JV2�>��[�ۉK��<��%q�W�)�T���y��40�	�iUe��\�U�ִl�l��<z���ן���Em�4w��|I��u��\�p�X�|���zI��\��Tǥ �[��5X�h�%5�𡽄���?����\��<YdK���������+��H풖V�{$�`��)����j��!�[ؑ̑���R����T���-b���
�a�|w�N)|�Ma�VBMMif�R�@տ�|[ུ�
��CB��g���݉����0CV�~rI8T���4�yͿ��#��xF��a2�u����0��B�yW�|�VDa�j&�.Kz��ȭ����a^D��Œ!)�e�ja{�2Q��
��=!�xqyl\��=:d|�re�C�^�vF�<6�� J��~O��j"
[����Y�\s
�f�F�)��,�P�FԠjVu.�����JMq��F���aQH�v��Z�!x�_2zh|��Df#��F���I��04N���0��A�[ę!�-��WS~O`E���6��.�� �
� o�n��Ab�����h����Ċ��N�����*S;���6��:ZH����.��ӏ����d���<�~[b �[ڕ��<O ՞�7#���l#�(�$��0�ep��3�oX��hb��5��nӭ;èE��鰓8���� ^�|w���H���=�L
1�4��EVTD�AVm>ɀ��!ri��+~�X(o�(��]O�j:=��6��J��������U2�h�SC�l3&�G���Gdb�xE�C��P�	G�b4�>+�H�h�p����0A�7���f1��؍�e��gg�̦���u?P6�ϻ߹�l�r|�Y�<���$�����pI��dc���Q�F�mrB�C깤D�]����稲*!���հ�DP�P�sx%p[{9��qMH7����W�~wG�T�F�.�ӯ�p����Dݮ�b���RM���q�E����s�����H�A���lg[����z������/&�t�����+)�#�I0K�c�*ie�������-���RSߎ�3X�-�D4l&�?����,
4�(ֵ
$5��;�s�)N�W�W�����ψ�Z{�I��_��5� ��8ھXE���3�
ԣ!�fK0C����)nim�"�&xZ3EAmPd)��N�rTQlg�	ƣ��bF�Sr��O@��(���BS}A!�Yʹ�Q�:+s�,Β��N��.��
_!*5�G9�_O�_�G`�^�� ]�'|��5�U�W��EE�y�;����Q�~�4l�xP�ە��,Wme��ƳW��M?G%nz�L��w�@��*���*�8j���dS�,�76�ʙ�$��!@��%�9����O��7+��G���C�.�&Z������#�̭�<����Y[j4��y�d�G��r!�
��F�����Jk-E�7)��W��|`��0ҁ"P�I;~I�VN�C�]�j`��#7[1��{�`Ga{�<8���l��&:����D������� ����0v����ex;ٸ�>t����g�����$��|qQpf3<�)̹����#�S̛0_P����������}q
)(AS��M-�5�Gz&1�E�����.�I|k�l�n��&ŕ��5���#���X]�a�"X�Z�1!�.E�@�eX@c�{@��]�V���z�ݣ8i�:�%g��J @7�_�.�$q��6�x?S7EP~��\(RQ�}���4���C�h��B��%�f	W��W����r�Њ jq�%���b��+<�[�����p���
�t��*�ue���Ӌj&���(9 ��X��?��s0j�(&E�i�h�ӥ%},�O͈l����+͔���z�0Ϫ���Q�#�!�/���z�50.�E���:�=b�o�d7���!�뼍
�+�T�HM����,�6p"���q�8	��<��h����8�c�%<1t~�,�c��7�$��P���Ɉ���i� �=K/{�+S����C�4��KԼ%j9z�$լ���k���Ǣ��A�b�oN�����Z%-j�
�R+��b>�E���.�Y>z2�����CΈJ�V��ڥ^3@�I�Τ,��FrfA~ P?ܢ~@Z�ה���ah|W���.=���	�� ��W�]^������N�LķQ�z!��v����r3����%�)^���ν���'*l�>�ks �lö�P5%"�^�2D��H}<��J?��*�ʠE�����V��.�t�q������fyy����D�3���9���H!W�����X��b��!�yvW?C��;���5���\��Sΐo�4�bEv��6��'��VÌeT�w��i���;����'�a�GͿ[���7��\fo6옺1uW�
}�'r��W��b�E�/
C�K`)��`v�Zkl�OCKZǆ�c�X��l�o��!ʮ�i���T��v\�BM�[�8[k;&e�}�1�/�(��꒡/m�y�k"Ry���+-g=��ZD*��#^�1��N�S��Y�Hm�W�&6S��+�қ�n`B[�4��0$���gd�.�un�0C�t�Lckӎ��v x�ʜ:tc�E�P�v�����-2'Yj�!���8�Y�	�9�k�N�S8��W~K��ݧ��D�%�����`�K�3��ev}��69sd_8��<eZ'�%,�����y�����*�V���r��0̥���lJj,�����G3n�管���C{$�FsvE .X���G)�k�?�@���Y��T1���ۦ{���%�����M����൏�֞W�����̭�a��˝K��G�s�����P-�B�2����:D��7��YQˡ5�9�H��v��u�Z�M�ۘC3��n�H>�}�o�L'2pGU��F��sr�އk[^G+J�����i��t:["�����+��k���2�u�~��?�|��۞����odM����i��!�J��������￧�N�9�z{o�_����o}���Q���<{S�.Σ6�i�� �X��O��c)E�l?��o��+"��"Z��m�c�a��!"���}��6��q6�a�T���h�Q�_T��'�}0�����B�J��4��~[��:���HFAE��aQ�tc���5Z�����|��mj�^��]��= ���S����`V";M�u�N�P:��:�9ٞ�|����U�����D�%߆��������M��E.z�@�npD���(�]��x:w���P@��/F1aEUe<H_�5,�Ծ!Tq���{������{�u��N��`)��uw/����`�.���� 9��S�����3W�@-T��P��E�@5h^��I����m#`������lOX���i&z��Ŋ���y��0L��glweW'Ot�|��)�y�*_���#�T�J.I��fg�A���pt�҃u�o�������`#� ێ!E�'�λ~�χ[���o�B���A�-r������Td-)!80�X}�n½��������OJ.������'5o�F��z��\���n�A�G���5�mw��>(�O!���Hnꩱ��iV��	�!��'�..MvO9�c��j.ࡉO�G��])��hCЁ�V8zd�U�C��$H2��w&�g�D�0U��O�������hݞ��6w�0~~�?��|�_��t��v�Z(�s�E��~�Râ�W�����N�`"�5���p�Q�����
ZQc��[k���{j$����""�|��}K�����~�A��+*�*H|�F��Ѫ8n�2���yV��y���H1
i��� 9��d:M��ؽʟT�9.��O�˨+Bz�6}%��t�������~�3�7/�AO�-�Ĉ�G)A�A�0L/�]>�4m�ɴH�4�4U德�@}=�}]���T1X�~I0)|7�������� �������UUې�o�)h?S�>��Vvog��`�Uw9�zu2������x�����60��4��'�����qB�-G��a�w�H���qy٘J�G.(<�1��G�qR_�  �B����~����P�d\���g�"S�)?�S�ٷ�9mҘuű��{�\6������tk�����̃k�=�]�6v�����>�}���U�D���7,�v�_V�RZ���V$:Y.ad9wax�|z�
���������J�������[-���=�9�s-����2��Y�YX⿸��W���։�.t����Ϋ�n��i��Z�=G &..�T��]t~�8|4���;|�blw�
�" �����`Ժ��M�&'r��������S�3ls/
)�^���c��݋���Di�_�>ZA��ĘE�e��7���)]�TI~�eP��=p;H�)4-u����Ĝ�����G�C%�P�Dv������U��&�D�<�]Y��Dk=w��9?z�tmJ{�[��9�`e��.��(�j#-�o�E�L9?.�M%� ���j/L�b�e_���Y��d�P��`�e�=������7�h21Q/���m�dV&f[nс���2���j��	�	��Q�B��]��-荒���Tɡ�T&���t�k�����p�W��`k9�d�4�j��)1���dO�_�N���P�&f�N����'���iqҥ�9����8��T��\K�~�ݗ�~�7� ���.������;�E3�C$���߅�ɕ��*=de���Ӊ�X�x߻�i�OY���\�08ǧ��Z-��m�Y�4�b�����2N#��X(laD�M���H�"vC�������E���{���>9��U�/���/���;��q�Ҡ�E��CN��APޖ�w%8�:<�j����%E�Y���g�zϛ��O4����D �+�X<�kG}ȸYN���Oj�ِ㳻�bcn�4w����WvɌR�ɘZ��n��*/E��AD�e���(]�����U�*FC�@-�p?�{N�?-�K�b�I�,reA�l8d�'>��+q|x�E?��[��r��a�k�k���q��|.��*��(�>��cj��i~��N�xy���V����/�?�|�S��y�Y�
�>3�����,�sr�Y��{?j����@�����Y�Y�z/��})h����0���_�+)��Y&�*�2���U�[��	�n��^�7��B z��t/@Re$]۰M�8���D4K�!(�ĵO(K,',*�#��8�9��T^����%٤_���&���jȌ�w�V�v�,iߠY]���-@V�j����9�)6�����x'X�=�}l�(�V;��|��Ç`�s��[m����t|V�J��:� �����?Nf�)�Ƴ/NH����<�OYC�S�G�=��0Je/�J��8���L���
�B��"N��q��YBL_1����"��ܥ)q%����V��kM+�w�վ���87����������Es2 Il�^b�j�>�j�d5��z���~�!��.]]>����7N�j�60��ฌkN/�)��<,���%��([:w�^�fm[�L�\kje��S^���BC�D�^�/�� ���TǠ>s�Ҩ�d���ì��aL����}
��'�ϭu��.n9lݍ'*)%����$�`�1�cՅd��@r6�pX6���&���A�����q�-f��5t����'��~���k�]��hԜ�{A�c�$ALҋ��/"�aJ�wu��� \�y��6��[���to+$�G?F����W��/�~;,b�Yr�x�\д'���:.�:'�/eN�½���U*l��<�{�E�|C/�Jf^�t��CzEu��������=��*���W��n�������s3Su��|�&夫6;;��@zH�qm��J��j�|��.qs�D{���=��ZVq��a�`���E�kv������ǜ���T�d�I�a?��f5��(��-
��]����jG����N�o��~Ҁ�����˃������8�N���̼���D-id@O��`_���mh^�
�7�7"%�{s&����;�粷|��g߅_mT ;��G�>� �&t �d��T�Q\v?�N�Έ��a��,��~h�HNR�t�T���P�W�
D3�zFC�=-4���|d	�x���=:���G_���\B�a���p([6�ۘ��U��ҢR�����h��\�F��s�b�������޹{���J�:����龊Xe~�S��E<O>N�i_Jwc���?xo��`�u�@Z�t�kŹPQ����Eؕ	���/���iS��1���>�I���|��>�T�:c�
����c�6�m,��T+�;f�|Ջ���H�(.D�dn�W�8o#�db����5x�м�~�"���y6]������<�wH��~9x~��(�t.�1�P�F����]��� ��oP3�MR��Շ�b�-�����WO���0��$�н�Ğf�8]O�(�w���C�a��B����4��b^h�D��R��s��K?��i��T[ox<� \Q����~���~9����kzc���'��S_���T�Z1�v#���&XU���Vj��`)�����C�$��2��!�EI��vO��������!�i�@N�������b���h@�Y!6�ƨ���T;����=��鄅L��aO�ZsZ1��&Au�[���k�^�-��8BK\5N5ҒLJ���H��gD��:��}�wo����#�x�{%D&�'�jEK룁9ꏑP�sA��t�bۍ<r��J�jN�rǯ���Qn��.T��0��n�Q)j��O~�,��fgͅ�~5��\�}ۧ���&�)���C�z4�Kӱ�B�T����+��D	��y����H��ї��|Q�Lc~���{-��Wf�&W�ިKj�׶�P������X�Pz뗳k�����ωҏ)�����[�Vg(maz}�hv�&�u�����"_D��B�&a�A����o�L9F���{c(B7�Ԗ\���׏TQ���}��W�d������ΔF�GU�VZz����
I�@�:�\@T���_^OR�ͱ����8��v��II�9齼���~��=�5|H��&����0?��{r!y�Q�&�+p���T�Ĝ�.�%iT�U+��R���>����d��ї���G����-�l'��f���W��d�4���L�����uO�X��Qm(ɉ�b済m�~���������Gwɩko���2?ƨ?�����
���[g��ج�g�j�'r��~��S ��gtA��.���?�V�Vڇ~�.�v?B����א��T�a�K�VD�����_�T�n߇>�g8B�����s2g�&2+��'6��I���	Zj�BD1Ap�p�����hi�f'N�����i�J��gӭ��)����K�$Y��Z�Aߓ�M��ɓ\�`��9�䣮t�H3��5�w�xaA�PiSP�^��Y����
o����Ѿf�'�c煢���o��E���g�ߣ��������է����&S��dm1�E��$�	@�E,�n�r�kA�8�����:��*�O�m�Wo�����k�H�uj����/p�f���<�Z���ʋ��݃Ϛ���1?2�/,u�b���{������d�T�K�y�6��nJ�&���ꞟ�ʩ�~�7C��BM�VHL��x<-��[B[�#�Tj���vA���<7V]�離�����.��L��3��W�z�v�c�qB_`�"���&'Sr|�H��ߺ�����K�|�ό�v�t�!`UB�A_r��l]����g���{9�K$�-u����J�a;��|!���1�??�ϓ��Zw�000���� �]�L^.ܻ�v0���	?4-�i�L��IKZ�CE�ȸBӂc�~W��$�h�s.l�-tbzZ�9{����V��x�V���c�`Vrl	�������hn"��â����l��F����}}����y,V��=f48"g�h�/��T�HX](�jHv����pUR��-��|:r;���!X�!��nS��'R#�޴7��9;��i��~�ѭ�d@CN�E���q��^��*�t���uu5�bZ�N��B%t>-���*�*
�Flֆ�)�����>GLX��y���6��s��K�\"Z��('����ȶY�`�66e���p(Y���ѷ�SO��Q�Ž>a{����t��c����X�F�]=4�&�B��r��$!o������M,ne�OßO��(�|3�-�tn�	�RER���I/�H��9�=�ra-��<O�<.'t�z�ݑv�}`u��F-�յ�����<.;<]�KN��7@��q��"1����\�,'.H5� 3@Z�Sv ����8��{������(�h��6�=Fy�K��;t��� ��3�N7�l��p�`��>��z_/�`5� f�+�������L�PaQ�&(��W����Ҡ5n��G�ӌ�v�(N��ޤce�g�Vi��6hM��Y|=����"FĿ?�!�)Fhѧ�i��B���Ĳ/�P};�kgs�փ{�
��;_��ՍFg��igq�c�q0�)w�!�x �����}��[{�����*U:�-��3���:yy�xx��w��/Od����|Q��F}W�|,=�R���Q��.?���O��lFַ5`偭mA��c<�����"�f{1���uv_����?v���'h��]��J|���˚|��N�����S>f~�5�/�J�,�Sy�l�!+WS��a,���6�
�ÿE���e�uO�g3D�Mx[S�Шpu��t� ��b�g5�B�9���qr���.�{��~]����C����c׃Y��&�b�����a^8ڜx��ǰ�V�i�$��/���h+��˟�ʇ��N���L}��!�����/�@���9$G'W��jƧ�V	��N�]�f�Z��+��`޴d4��B��� /YN�P��ݚn)t~<�ߑo�T�6 �W¬�(�	����V���BC��/��$].k�k��;Ό&:?���NB-��˳���-����)n����ޡRs�\˺j�[)O�8� r�兆2�����"R��ӯ�`?.��~����`K���^�鱘��k���q�����l��`ؓ��������z��	��b����[�U�}U�K�fǸE�Z~l:l|k��O�e,�
Q�ܔ��w�^�{JFt9+w]\���Ԙ����잩�G�(���/��������#���Zi�RGg��$�豆|����$Upbz���{�ǃ
��w[?�����H���_����.n�T�"T�w��ˎ9�~�\+�*���0�]OD���e��'|�쮹����m�q�RX���p�@넧��N�ɬ'ḨjV�ߣ��燆������"�_����0 ���@����V��� N�ƠQ=�h���_f.Γ=��%��}0:\��8Cńc	����K,���U�?N���<�w� 3k�3cҶd��%�x�ÖP��)�f�T�D����@3���1��}���X�!{_x���1��,��қ�N"�殇�7��:֚;X��
]�t��X�;_2�QvϞ�O_êа۰���e���%���Uk�����n
X#��{!a�? ��zG�����{���E�\9L�1b�8&sy#�����p�:	R�b8^���x��K�������Q0L��t�\��~b�U�;���l�A1�W��B�Cfj:�����[���;���¯�$�������+�N��~c8m�|�HYX^�I:�
�rE��+�??͢bl�%���'��wb^��%�M�%7�,�p�.�(��� �Ze
&��ֱ�U��zHj�⒔SxG������s��x�}n�	���76d"�0����d|ւ��t��e|�>�-��<f�2V/�����l�q ؅�ߗ�7?iꊚ̳xT9(Mʭ�k]�XRr������Z�"�@f䜴���{=���z��mW��D\׈��a�����H���h�QeL�)b&����nxy"���O{T���Y��]�V�׋�Ttp=��$b���r�3�R�y����F������<	^v�Ɛ�އU\ӟ�`,� ���%|���Qf��;�`�۝�z��b��0��:[��B���+��m�u�A�Ja]{d�Gc	�_�=M^�j����[&h�달�uX���4��?Mگ/f{t*O�Y4�|<���*���l
�&�©^����#8
S��w����������8�t�;XÍ�U��{f�.SB��j�
�tg�G���rc*߀<S��w���Yw�cl���[�A�ؤ�v*�vȴ&��^Z�j�2J�26յw�5��J� �]?;�_�Xv\�2��N�h���ݥ���*����A�vȪ����|Itn*i����q����>t�dғ-��p0��0��ۘ�e[W��l�8�5��C#q8�i���89<b2국D�M�Q$h,gt����hE�e��h���ɯ��_�w1.�	��+bƐ�G��� �6�ǧC�CzU�U�ܘ ��f��)�K�l�V7`�S�����5�-�LMcچ�e'��k�[�N�����c�cz�!'Qt�5��3��g�)����#�˖7���@|P2�eU�QNX�k4'̤zp3,�����Y8	#�fY'Z��v�%@�0\�=��h+��m�&\�NĬ�n�
_k��Au3b��?�ˍƊ�8֐t#;V	�����q�g���j�=	��ͼ�Hޚ�B���ـf��97V��i�����F�qߜ�370!.�OWT����j�2ڐ�����ɦ2+Se%x�p�P��� ��\6���>��T��Le���q7�,���)>��9P��t-/5>�>�4��ŵ�̣ۭeH�+�!N����U�'[��B�q2���5�K�x] h=I"�fXy�{)�f�5GԠ-՜���`�B�D��d� �3T���m�,k&M͜�����0UL��_c׿�ӅK�ٯ�-$q���N�S=K�ڵ��/ݬ;�a���畴qts�{El��TGs�\&LBF���X�����-���)G��܉3%a�厍��j�x�43���ze-Q���sN`�|�g�E7�#��I��u�d����F64�Q�o�W�3��QQB�.�Č�$@O���q�����bpT<����������V�`�uF�k��Шԣ	��!��&f]��`���O�_TA&��-L�h��8���!�i����wC�Hp�{�D�mOkF@^� �G���4=r�-:�[�˛�M|����s��$�1}��Aj�`M�o����ze&r)yx����v��]�p=�e$r@cB�b)I�!��I��Yvi�S�6<�Q})<���zk�s�?�/�oh��6ǫ�u�"�#�uu*	���r���x�x�b|n�b�N��p��w��-���;R4�e�o�g�Õs������ŕX)-W����ڛ�?���IC}�51wH�=��HU�<a���"+������W�VW�N�uA$�ޛ���[Q�'�����m	<Čgt�"�1�BhR�Z�F��-����j�<����p�(�
��u*�^�{ċ^AP4��fw� �=����A�)��Ҳ��*���O	7I���
.�J��.��T�3p�ŁΗP�c��澠t��}@v���o�ɋl��B�E�����,�r�)�'�'�n'��S��y��38pj��m�R�o?p���v�L$U�z�{E@�@:V�$������(�X
�K�
2���q���Dژi�:������}���r��"QyM���W��S���p�����Y���F(>(�c��D�?�	k�v��2Y.�^*�}th�)�D����2���pή�2E��5d����W�Q�N�	�wC��F��º�b&��(By�J�1q��<��4;�nബz7��Ni�/t�Մ��ָ�X
a�;s���2���x�g�����ZJז+�ɄtN!��e�ذ���|jZ�@6��Z��I�PN,9���fR1}����8�E��)R�N��#:�4�\r�ר��Q%)!Yk�J:AzX7Ӻ]�Y�@}K��Ta�?����*!��KVv�Y�YKL��Wг��,2t���;28�05E9ʡ!�����+��#%���C�i3��1`�X=w��8�G���X,I!& Oܱʑ���+�R��T�ꎠ��	-��b硭�z�s�}�I��l���5����BX���]v��w���ԏ��!8a���'@��N�9���n��+#RK�:�gР�NbD���:���&�\/o�=�Z���G}���{]|�_L��ԇ
����D�Sx����W���1����xO,Ǜ0š�Q$�? @뿪���Ś)q3d1T��@�K�2:m/�.�r���d�|��=�.�!r�Ήp#�j�H]MNϖ������B�3�i��b^T���r�Ǫ�;��2�m�Te)�;b:�ؔ��܈�ue�FK��9#o�T��nC�:�H�4�9�!������b���J�"W7�5Twn�^-��͔���
m�M8�ʲ3t�8)mǇ�T�72�if�\c1u�n�w|Qfn�TIB�TrK�#�h��Ǡ���R�=��U8w"Q�* ��XH����$$�{���A
��|ȵAW�I����e�W�K��ρ.��	�7Wܒ0E�=P�:C1��X�
�7���!�0T��%Z]c"eC����:��a;��^�K�M����]�aXR�L�[��78�>���w'Q���*�U	ո�^�+*a�,T\�&��,�Y#�7�2]Mݶ�ާ��UR�c���H޿���8Ҭ�c*�4���	�q;�+���F��������7c��fsyD݁�M3�|�R+(�nm��cXVL�k��Y_�T7f�rL����i�
mc���G�a��	�D
R��l,=.a,�2�9פ��a�ed�E��FV?aX:%����-FG=�8Q�c(����p	�֨���k�8���$�p]���
���M��*7��jA&�p|��T�\C�4u>���q��$QjS�a�y�������@��1Rn��S�aR�O�^�����s�����3P��ⓩ���춹�ʯ�Wuv�R,pR����H�2ajk�D�W*�����D���^u�ҿS��M�.��wc��W��Z��+�)�ߤB�ҡ_���&���ȥ*AF�f�N��o�j=;5����aޱ�׆
�]%�UBˈĹ�֠��*��r�g)�I6���qX_1{!�Y3i�Cl]'R��*���LŸ���`��a�!J���ej�F:׆23V	:U�~�:�*���]!ŵ�a��^�Rảf�Y��j"����l�pMV�Zp�<�.�y��k����%��h}�T*��i%mT� ��vnڄ��L}�^:����g&T�OF���%W4�a�6���M	;Vo2�%�B�Sc�K�U}p�%
����(��&7�꩎�-b$�
�Ljk8��*�k	~�響�}�#WOg<�d�?��B*p��GAV�V��ޙ5c��?��Z��a���J����f����U�����z,͎_���0Ե+Eƈ\s�ᕮE+���uf.}D���Hʾ����=_��Z�d�yY��?gBeU����1��$Q��>2��j7�u]D7��V��[���q�-�yI�ew�N�Ɇ��!\��s6�dV��0J����[ffEP��3@3�1���[�I*�.�W��gK�F:��U�����ܒ�0����(��*U|� �k�+�L,�	|�Gjßa([����6 �:������0��l6ތXxl�
��r3�H�.̟	U/1����A�UCj]�X0T;L� ���`�Z�n"�~�LU�R|�I�ѵ#w���˖3�@�92'�ؤ2f���J�U\��lY��*S���A�^���TG\c����	,6d��,�P+�x=4����� &j%pq���t�/��T��_]hfU�WW��d|����87C$���n�a��PR�k71]��
Q���
�D�J#6��2d�����Q�0��4�Ȑyku��+��Hl�bIk[k���Qk�߅c�@-�Y� B:|���\����s�ʡ�W�jQ՞��Nn��)I�^����RϤ����{�0�\�{�!ZI�+6�A������{��Y��H��Pm໇���*��I�Y����f�,	���2ƥ��2��>����ԛ0�J3��J}S�e4avC��گ���ߕ�2�S ����9�;�]���ʧg��*�Y3�ֵ��W�%+KP��K�w��Wt%�kz�8vnMS`%3=\,�L<�-n��Dj�$�WQ+�ٜ�,	�_C�ʾ�=R"�B�N?礥<��Z���wrXD�ۼFw��g�~���ZۇJd3Y�:(����2R�z�;��@��((٩�ʃAOIC)��ٱI�1P#c�	q�ן]�B_U���O��,M��{����@!���]�#^� �G�7rf�3��e\�@1#�)�T6�l,Y�qs2����^E\υ��u8&{�Jx�-�	��,O�F�^�A��17���L$�����C�&���?�8|^%��q�@_WB��0�*�Q�@����{`q~��j^�h�0��vƙSUV��0/��rofQ"��%h��TަJAiI��Ū��1M��J��A�Cz�(�O1�( Z2��1������L<��1���И9,W�஢ utU6e��g5��:7����$�ĶX���Ճh�j�U�ϻ��1qh=L�Տܪ�ġ��F��֖��C���˜��T!X���hV)x���"Z�]k�]���h*�M>k��������c�'�����)��	
N��Kdj��>k��5��^ψ?��ͮ�y͸^Ɏj��.�l�$�1�㵾��c\v���6'���Xq��B`�D�1��A�r�A��ȏI�}��W̕���UU�8�?	h�J���k,O�bŮ�ʃm���j#�0�0��9Ώ�Ŗ��"dq|Ǭ�a��Ư�:�ps�9�,������=N`g6�iV��/�>M~��hIc���*�\K�D�g��!��� �V�)�}Lm �5���3rz��`��3XN��Mj=R"�������SČ�j$�-���?�NS[�H�g����W�a���G�������	\�$���P�+ү���B��D�7�z�P�MǓ��e'M}I���
����X8�f]���z#�~H�={�ޛ5nH$b\�C�{���0j���1��bR(&ц[Az���ژ��n5�Qߓ�:�?�Z���k�H�gߟ��t>�t����YT+��HK��ހ�B�.��Q葎U&���i/�b)H[�MJ���T�΀2@��2Ie�.����	%�Zz`��#lpr�DB�Yg��nwE��:Zte�wZ���/Gf��x�jP0�f�n���76n�"QQX�r��Jc��UF�6&I^���%�|կ"e]�,��Z�6�TI���r���?��3�0�K��X}="�A�-�-46�VO֑�K8�R�$�<&��}�>��@�\&� ��I�2�e�_����cbbJ���i.%7�S|��2���b�=��D���O=�m��>��}�!`u�R��|�Ks��)�</�r�����ѡ����eFJ��-�SϮ��b��{��-�=Z�3�y�:֡Σ�Sayp���� �C4hhƠ^_k��~���*�1d&���&�2��C�TW�mT�^7>�|�D��B\��F��.�Y��r�7��/��N�g����*�UC�&��1���n�H���M4����&&4�v)A�6'��T@�6�r��TB�}Q������p��!f>��R�1����o���}��f��"=u�(���L���%���/�=w�m�h�Ԉ�`ˮ�zM��:��1��o�>���ӈ�t�	�y�$�;t��ߍ���w��~G2�L��8o�$�Ԋ�h�)WΙp�1��$��e��ex�J/6"���ʢ�4���.-	�5́l�,���Mh��M�| �4��T�$o.�.����v �����s��yT�)t8n"������G���'U�VŠ5G�A��K�qL��x�]X��03s�S��VC����tۈZ�t�.���Ǡ�HC���a�;�hG�~�m-z�H�9♨�Z��J���s�؋O#�S,�p�4���������=,��6��;�P�Z�:?����$�E���D��ѸR���\�N[������.16N_gF�jdVY;�H����uB���<OL�9�T$l!_��A�&KTNS���O͐�2 ��蘍U�/���5��=$�bNR &k���2���Qk����l8�W�ҙ��ߛ�_��(ߟ����Dj{��ٸ��C�g#��m)<%�]�	�lcb(�7-��0}�K�Խk�	�V����B�f>����2��RR�v	NdɹBÌ�j��]�]�����v���p��֓31X���?2{кz�+sg�]�ν����0�m�G��G?���u�(�����IƐ�i\�;�i�lV���m�%�A*��v�B%��T�j;���̅�5�p��Y�V	�|w_I9���Aq�Q�*Y�Kꁇ�│�v^Ar��N�<��"�E��6��;\���t:��}��1�:��E(�Q �����h�hü>�0sդ
&�1@FER��H܊j!ؙf+��i!I�>���L� �i-�O�btt��UXo�La���k� �������\�6����7���Bc�<����[o��e�XBݕ�{�P���ʥ�����F*y����1�>1�Hi
�K��R�Őtu>T|`{��0N
��|�v/]a螗��c8�ܐżʋ�<�2��Gʘ�3�a��ÙI�L
���{�X�B�O���9d��-W>��3�I}˻,*3���e�тx5�ݛh���^� 2X�9Q��:�LO*B�}'*��/Y�^�e!�<�������P�3�L�Щ��Q���=Cp�CԎ�co����d0?�R�A��� Z��EN�C�jͤL��TQ��/�,��������Q� ��V��?F���/�����,�'�1�I"5�p�ҁmA�g�13�&Ɏ{��y�l��ز����"W���K��}�Q��bg�R��v���h��D�\;!'�5:��G�vE�{lR38i�u�����2�r���'$1Z\ۨ(u��
Ӑ�Iprr�j+�A}Bl{�����(�F��������旟h�.��J�E�MKh��W�ѐ�Q7�]��J�y9
v)��������	D�n��8+��D|���E��)��c�O�쓺V41���*T����[$y8[�e�xq��H?Q��f���PX�`r�,w��ڸ|�����6�p��9)8�M��m.��Ip��Y%FAh!��y_ܕ&��G'2�AH�3g~L�!2	Y������%��U�R�9i�d���P�Ab��A�=Js��(\������
�h��mr��&�Xɕ;6T�M���=�ȼ)����r]k���C�(�(�$g&�X��!<_��4���2Gt����H��@@�,$�ÕN���jZ5h[\��PnU����!Icf,��Ô-�9A,�:�x��5)$���˕'���K
���<��*���qx�Sf ���w��?����*n�9�i�_�����o��q���x��0;W@ed�v�׳0=^D�@Ir�h:h�����c�1 ]�#�W��Tݱ�J+������	z�@�ֽ�..+�$�c�KuT�N ��1nQR�9�m�.w�6U�N�b��A���0�p	2d�TU�[�h!�h����`�fb���,4�.���'��~_վ,%$� E��w\�����`���hs�t0<BFyF/`T�ь	��<fSEr�i�T�`ڜ�k�)Ӂ�=Q��@.�͠3{&!)z�J�"���=K4���&�E��a8 F�ފ��0:RD�PM}tDr,��H���bҡ�cf�wI�]^����E#�:ĸ�4'�����\��O*��\,�Эs��lE7͖��jKڴ
�2%�S��U5=�s��TA�$r�ȏ��*IB`:�pYgwLEHQ��擬���P��6��E�l�Y��|�����u�UUD^�=m�Ȭ#��>�,x^��D��0Q�zbF�b���X�Ha��pYS�EUFq�I���$%L��,x��p��%�����h$�s$͞UBAC�*���UTB#���r������ݛE[v�a��3�s�g��������eQ��"��-E�W�V�W�d%/^+���<d9ɣ�N,ْ"3E�M��ř 14z��w�|�R�U�{�sn7  %zSPw�{���������*�t��1��(�s���#�K�?�"�h_�xw�"m\�>���Ev�#j���׻E=vۇ����w�7�Tm�fb��67�鯽@/���ӻM����yb�V�%���SokD��E���m~�](������|�ۼe�^���Ke �Ga������i_U���٢��%��s��cmSF��G�4�	Q)��M)�2qr�%C�T�R>��v�-z�z�$8��P�X�Hi��e,�r���_��Z���3�ϭ�����S��(����p=��`Vm:��C����qH$w�p�$mܾN�`��5Kci\4�4s���G�:G{`!P��|�t�ۿM��mZZ9���]^�ٔ���1���)*w���&����׮�djE��Hk=��m��Ʌ�Y��#����[0�@��d����'�Ń���Hrv���P�7�Q-��2"��5M�)폌@�.��Tt�+��W}	�$���ҭ�f/�#�;�C}��ǏJ��Pc�(!r�4y�{()L�(����ΐ���L �����6)���6�Gąe>���b���w	5`$#���8�'-���̥�����S�T;D�*��+��y��4�B1 ��]>��.��G�?���x��{�h�S]�6o�D�{��ghaq�v�y�q�)hn�"+��Q���1�`=j�t���K�?�t��r�v�h�4�����)��������TbwF"�9���mmt9�X����6K��tf^Bֱl~U����'퐍V�a��6b�{���<�(�֟��V��Ѹ�M��f�&�^d�:�C�w�j�t��� �&�1�

�{�9l��*e#l�I.JM�ْ��xj܅\"�8%��LZ����M�۸A%�H����ᐫVcC���R���<�b̞�!�A�11�vg�6�G��m�;�Og�����
��}���Z]�B�n�{'��ҥ
~5�$j�%�1�� �F�$�'RF/���-�y��,8��;�մ`�Bu*AVX�w�'�0ACP��EFVJ8#�ۄ���X)��%�ȋ��jRS���=�*{�=$�� �>*XJ�B?H��,�d \m������M��׌��>#X�o��*"皃���e��2��-�[3�q���ոJbr�ԗx���	Q��o<���zJ��a�ׂ~��HF�ү0�b�a��,9/�,�y��� �0@"���u��\g�Ve�����o�=�m����=N�}����_�*=�oC��Qi���NNG��
/!�����ԥ�G8+�lu6(j�̅t�FJ���9:����[���v�2D"������^O92�#Rh ��M�h�:��H'F:]<��Z�2���X�J����i�K�Iu+^�}j���d
��-Ѐ�~l��%>y��]<�����9�xD�V�q�T�>�rܥ�?���%j�8C�c9��=�dp��X+ȕ�^z�hn��������o��~�^z����6-�� J��<�C�Z�<���-jq�P*W
@���N]t9-Mf�,2��t��Dbhy�T9�O���E�
���� �l1n�t���8�|u�NV��F�O�3,=)���[jKY�%�*Q�h|�+����e���԰�44�[/�j�xʫ��*kS�i0�tz5�5���ךQ?E��AjUu��c?&`�", ~���;�
���3�̸� O�+g�աc%�^9()��(���VϢ�����\�5	N�����滨�+Z�y`"�S�)��Z�����d̓�ߧ��6mn��~ϣ�~���}���q�#��.�S�2	e����A8��4�`	�;�@��V9�8�F��������O���Ơ�@���#%Z\�5��J6�.Z%�8�Y��(�&�'�o�*PUI{m̋p��؍JjI��$^ܴB��[���Use�_��mD!��B�����3���+3�a�����`e'��AVb���i>l�ջE_��?�o��7�W���_Ze�����ga��!�W���Sq��-�Ԛ|ܟg1�>Gh=�bUE�<e�������5�"�&�1�>n��x�T��!�NTO;�����]d�����V��58��8_��(ֻ�ɞ'�0� �ȓj���sȦGſ0�ax�%�g�=P���G�g(��ܯ�Ir0B(blC�7�c����~�zZ��]�R�32^^!�����i�1I�'9�
������PQ��CPP~~�@֞�L1�������2��?���鵋D�]���HנY�M'��2 ����޾�N����Hυ��#�����{���-�_������F�A/3����s�����6ـ�c�E���{@����|�	F��s
�����[�d��|��`\\��
�i�{�~U5���Q��bM�T`l��V� �.ě���^����[�dO:�w�I9ImI�	�a����,Ǔx���BL���k�����Z<��8s�5�����NOɑ����,�,����`L��3F����y���
�S0�K*r�d|���R�9��f)c]�!��J����Խ^�S�N!Wd�"K��	�`�r#��Us*�qY�J��q�p���#�@3/ g�{�XЋ d�lΈ�e�OG2��ʷJ�*|������}u�[⩇�5C���@H��Z�K���}�l_Z҃\�2��8�,��ɘct�"��<uz�Z�m��n����Y�����:q�8jp�,R2��A,��E�jb �ȴ+x�'�$�{��	�<��&�M	��j
�&��?Qv�+'w�8�+m#;+���Kz���e~��p,�JM�'ኁ2݈b<\�@%�(���4IC��ll�|��=������J������,����00^��44E�
�ք��1��I��Y�Y����4����L&צ��ϖ��촒J����7U�Ѳuy�X�nt���9�]dH�rt���O���bρ�l��}Q3C��pu=4��S���KF�3�`�3ͳz*���|���}c�xe�
G"u���
����Ce�y�&͋J��`��`�C����"��\��X����ԣp�*a�8~ �I~6Ƙ1�vwwh�G��G��:-��w�:���G!09-��:y�DU�&n�~�Ξ�@{�Щ����V�Q_���1����<�v%�*��w}���@"(9�S^�:wʺE�z:Y�Lh�ad��𒂁S`�R��8��!֮�Ѝ��OU=)_.�����i�. ,�'��s�*���0���}x�y�$	S+Q��"u�jt�ɳTi�I\���Wiy�E��)``�B��ԨՐ�#��P;�	m<���T��3�v���A$]xn?8}&��_=�i�$6wS/%W��5J}B��E��E�T�q"��a���)�}M��0��P�MS� ��QN�Bw���&#T�]����%��d���0�6��xO�B�����
!~�$'=G/�6��* J�إ�:͜ ;D�o�I= �r�H�.g��L`~$�ɩ���	j���w�UpQ�P�e��4e�no��?y��o>�'��T}����賓yL�OA8q?�[7n���{ϟ�W�Wh�U>Q��c{U����-'F��hJl��xN=/�׽$��reiq{!��9/<�I8��"��UVe����V[��w5&��&+z6Si5U��-����X�H6K+XG�k���n�v������w�L��|�]�.}�������SВE�E�A�c)��p }DZh#t�4���kiI��u���
�ĕ�Sn���siII*�b԰Ƚ��;D^��(ʎ���#��.!�!�z�H��Y������`����m��lj�"{����/5J���K-7��<�R�,��a��'�}�H�h����|r}@'�[�����Ʀ~/��IIgvI�d��J�}}~-�OM��Fĳv��b9��z���qj��X�/�q��]�Q�ݽ=����{�_J���!�f�P�{��:[��_~�V�f(.K���?���W*%����~�j^��aH#�t$6!:2��Wq�j+��\��J��+lH/)�$�N�XS}�?�t�x���a1�� �7��5�iH�N��H��N~�NƉ3�n�.�����,��/ˠ�i~�I�M���eϳ4SkPTR
�h`��D�F0�U�@2䣨O�� �No2�]Hd4.ķ�3H9�3(%Ք^��K�!AA�kT����Q�<<�OX�X�v-��g���čGjd	�ǁ���QIV�/O�D������Da�f��ϼ��<�e�
F�����j�e�����@ev�8��l<V/90F��.2/!� ț s�d�U����)��XDUM�|n�XƄ`${^d^
:������gO������
Tn�[�Z�����[����M�׎�$\�פ /�fJ�R����ԏG4;���߿D�����O<̫����볫5�P$Ģ�Pv��l�m��Kj�ڂE�S}�;�a�9��'� ��j����^��;�y�.���G_g�QD�'t��v��M�0懝�ӑ�e�|���6�0�gw�vi�6Km��:Q���z̞���g�g�$Ք`���W����ધiM�n�5h�A`$?�wK����N� 
J8�pZ&�����Q�Q,'$"ǒ�S�>��D�`�G�o�)V��;�*�G8i��c�>��~)d��)1�)g����k(�`��i��1�v6uy� ��h���S�x�Y��j��S�<ߌ��B�V�N��_�9(8,��%���Υn����3��<���ܵ{ ����&Z#>��2�3�uz��u�ͭ����0}h��O���̯��4ÞA̱p�݆��`�>p�Z�����-60k����~M��%���Hq�F�1��#;lҲ� 5�%50��g8�ssI�s{(��ْPs����1l��Ir<G"�[��	ԟ�@n!�X�~Ow��a>�a�A��'�ě��ZAF�Go҄�!}�2?�q$�rp���X�AQ���R�#Tk�:�͵�^�'�)Mh�^�C�1(V ��2��擩s30���1T�cd��SPR��bf�x�xh	�͗�4�HOb������%Aj�O�g��֐�]�ܸJG2��g�d�������FI�W�2��"C��k�蕸�xq��|��Ƶ�C��x��_�=X�hް_=5�e����zf�ū��.`���1b%�0�!<E�ޘxq�K� �6���0��Q1}�֝�T�P�Ër�G���>C��c�!�Vݴ�6C�y:�]viC�f��r����O����ah֍O=��(�/ŭz�]3e
�].�Fވz�o��`����x��A/�05�������U�Q�D��5�\v��
Ƨ�k�^��6iQB��C[=��3�4fbƹ�g"�슲+���R6�P֍�"^�|p��ݳ� �؄·��v.ˆ���V��u:�d�|Ф/&j�q�%���ƺ1��L���:��ÏT�q"�S'��N^9�m����@�P�(�6b�gq;%MF.Y�(O�7�d�Q�����g�6�&��F*U#�Y-��02�ًtB���$���N �ϿW��i�Ҳ1Z_�r�.R�>0��ť(�Ʊ�u��ߠK�vI�6�+p,u�O�M�:%Z�"���\�ם9y���/Ȟ�cOL.mz���Ş��B��[?R��]wȅQb�?r�4u�g�;���ߟ����(���h�S_�N]�������7!����ٚM�_\��. eEd�M,٪!J��&>O|�P 7%���F�V��~�8]m=�@E���:9N�j�C���g�*��/��X������l�6��J5��7"A�< �,Hcv��,z�$D�iN����	�j'��k:ѥ�5e�n�6�q@�^���5�q�w'���)M�LM�
�*Ǥ��ylϔ ��>`얡A�!0=T���Q/V��{F�{Y3Md)\ߍ)S�	��<u8�ж�~��K��3����*��U���i��(j#E"V�C`��_�Օ5��@	ʕ��$�7�5wyGN�;_.&�t ���o�*��X����4���]���r��-:��DK��x��I:8hS�RCJ����O�[�K�T27��_N� �]��)߿T� t�k����&Ȟ]�r�T-Z�f�YV����V4Ҙg ���*{=��@DR�^�j�]>�J�uc�x#<U\C;�%�M|�}�J:Ԍ_�8�1��>+�LI{kТ��l�f?I�K��.�fB.��Է�[�J�WĂ����#4�]����*���K�B�y��v��<"8{�u*%�L+��g�B�[�����쌨���hphJ+j�*I�'E�ŝ=��-M,����r`!b�����Jv��8w�Ҍ��?�[��,�xgO��w�����M'?�N���f���t:ܚ����,t(�զR�=��)�3���u���α�PC_!�I=C��i��j�܁9������9$�1p���ޝX����{�� ��7�@��;Ue!�:C�&p򩈌�pp*=:��O,,)�*�hS^��T2��v���M4KA��|��-�I_�a�la��J7�=Ӗp�g(�e����	~���&AMMA�D-Ou�H��j��Nh��W� �f*�F]��z��:~�9������^����	1�/"YHbU;�67�iqi�~�.:Apc���p��-n�+qC
�VW봰V���9���l �T��Q������{GN�7��&:َK�q/�NWƼ|�G|{E�Tf3������.U4;W�4�H����@��F�5�*,�E"؄���̧�6'�Q�K9.���[Y�����)I����+gV�%�_���4�����$CUJ���}�����9%&g<?rU����	bm����H�s��fL����㼇�dY����{N�W�d��u���e,J6�ƽ��I��e!C@.�*xKj�u~e��D�^.��� ~	�R- t5#��)�2+���]���qDB�@�46��p�S��kЙ���j�7��u�w>iv�m����TG�إ��y�ݣa:�W_{����2�K��X�����4���l�L�pw��k吨�9-��R�Ҿ9�,.���������I�����Ig�65D��ϐSWz=��	�~-�4[���u�p46)=�&*a�J%M�n�Nd�� ]���r��i�Y�)�NWY3��ȳ�Z��םĨ\tYc2�Q��R=����IPP$=��D�n��"�4�̥��FS�ˑ��qa�����}��0�p[h��V�%س&΋�����B6\��#M��12�0���i_j�D���Z 7SE�b�[��+f�XK�y������
ͫ"�>��_�k֞M�*��OD�B�?#u[D`s���N�^��A��o��vL��Y��(�����#*e�:8$^�)����K	!J�ס�E�!�־Cq���P���k�O�~�N�}�"U+�����LU��>I�P����ѭ�Mxm�z�Nd� ��D-�/ى(�4���V�c��u�$9ME^���0T�Ps�1�c=`2���<�[��vb��2�
�8�o�Z���
*Je�dS#x#��������M���88IR]P1t�z�YcbEgD�+�ӑ��%��	{�[K���4��]�o��:��C�"�<EƦ5o��TO3C�9a�y�!�>��$!#�i�ixq�s:R-�֪M�q��#���)��2
^zV3ʩ��;ʃ����׾Ǟ�Kt�;�Fc�cZ��\w��M���=d;���8���[���kX\�->ͺ]�i���X��������e�ȸ�8 ����R76XSi���6�!3v¿����.�.����s+R��$o
LȾ7�;eS���o��g����Қ͹�volR��7���t�(T�ֵm:u�4-�.��=>�y��U���%E>�|����5��� K�^�y�R�'�����UU�9v�-���^�%�HK:��>�F�p���9�L�R_E��ھ�R�pK��Hė+3�����R`nȐ(��y92wq:��{�G��aSZg��:�=B:Ӳ��|%�++����K�P凪�		�i�K(�j \(�����(��[Rv�x~����J����c���B=z���|5&C���G�����ax�:�����K��եy��O|����N�;��(�5���`!�H:i*����D�TK�P��XDYc�<�Wy�(�C!�] X�*��݁H�|71�jӰ?��w�ӣ[���ݺ�A��7�<�s���3��EQ)v��s��BS�ġ�P�ԟ�^6�(�!D�0Ӑw'�
L=�2}�����	���l�X_�*Q�@7����.���$����c�a[�;*LVǑ�$F��2����c�^ql��#��ֻTkT ;��ʾ̂����O=�(R� ��i�S��r�3��3� ��f�FU�;0�*/}+;���%?o23� n�y�0�?i�(��Dh���q(\Bv��Ҭ��S�ӥ_���l�΋��q�tf MI#^�}�-/2Qu�!}D�I����@+�P ��o��e��4��c���r�ֲ w��7�b��onh�l(�>&8Ұ���]4�A�o���{�{t��.�\}��[��Hm&�=���x�-J�k��d��-0д�~���&7�߳�]�����g��&�R54�I����G(#v�U�&�;�#7qx4�S�RB�#y��N�4����fɬ�:���#�n�6O&Hms�)���2,0i�YB�4�1�ϱ�������ea�S_٣T%W�I����e_�a�~�+SOQ|�v0T�|ˤ8�K�z��zobM:��N�!��`H�a��k�LXx�f���a�b��Wڴ�J@�eq�<=��Ef[�"�f��1�'�}�G��kt����t׳���~�Q�ǌD^����r'��+�C;yM�b�b���iΣ�u	�A�6C��U��u����DA�ĕj �頤�1"m�l(
��`���V�'�PBBK��1ʤٵz��9��Iiʉ��ظU�Tb4vL��xF}�5����F�}֓e�0�ٿ�vBW�)n(FGx��6�r)�X8�]��S3�����Ja��l�2>��L�S`z���y���� #]���֋��O�c�5����*2��K��
5�4�O��(��X�t�a�c�����eцe��H�I��ǥ�s�4X;�/}���	nekƇ�Sdݦ=���ɜ�)������v�'�T1��XZ�0(��.-�I'���N3��$�Pѹ��N��o"LcŐ����ם��B�Qv鮻��F$3��g��h��q��!�A�½!]����s���j�����5�2�v��l6��[��kA|	Yv��Ҳ�Q�^��iOp�}�Y��M	��x4�w֤K��U�
���ρ�D ���U�%0y{,`֖k�#Qڮ���H8,�/hʛ�O˕ Ս�����(s�S�N,k`-�p����fw������t��t?4�w�F�j�y�!(��e��aZ�����Nc#P?G���Z��|�)R'W(�����<�3y��A�6IͣI���R/3*�-���4S�t��*�n޺Ii�&�(����T�U��+4�-%(Gp�Ő����(JA�oL%O�E�'#��+�� ��	����3|����g��f��L��{��̵��,�~7�n��(�V��)�^g^�B�	�Z�i����������z�ܐ���`��ꒌ�$7�8��'Yz���O-�6���f�����T_@�
�l5�R�;���-׃�����GOC�L���QԦэ���e�"��d��O��������pd�vt}*�|�k�p�T��ss9?#HA&�>�K��Uq$8�k���phAY��u��&�/˪Y���$��3U�6-���yË��O=�Z"N3�Q����S%P}Ji:�c�p�{H�;�ؓ����.���=ԛ ��WK�D;������;5��gm7i�r޾���7ry0��SZ=q��F���*�����1o>)�ړS�cc��DH�n�a[��+6���#j%M�N���>�Y(G&SU��(�%�lS�^~�Jؾa�	�dE�u�pM��u�ԷjO�@�q�d]j,�l�}�n�"S�� 	@�����\�IXOW������-Q�4�>R�N��Y��_>ט�T1	߁F��P�<�3��L�!p��ϓg�VCjrw�C�*]��A�����ݧ��h6D=�=�g�'IR�"?{����,">R2Yx�DՇ����ѓO�4�v�"}����^�����R�S�p�ɓ(����>N�|A�K�Y����ZLYl�����zY*�����1d-~��K\�s���_�h����'�`��������4�uz�{��H��s����1�2�$��������)l�>!�ĩ���@+%E�?D��Sud��EY��Elt�h�:/�����	��1�>��啈���;�t�{"0a���Fj���f@��u��SI��
�44 �#������?z���l�&�f,T@S���U���ħ&�&&�&FjB��f�o�vG9W���}慘���8q|�$�_xy�p(���-�L@��K�nn���-�sO�"������ ���pb��ޠ^��O-�$u���*0�c�xI>i�j�̨���xV�n�9!?_�#<�t�u�������i7н?{����~����%,r����u��o� �t��-��ܤ�/�kԨ���Z�fc���{*8��K���T��<K�!!���rP�72�����4��Þ���7���d�׬/����`�ք(�pd�Ĩ���<���K��8�"���?�MŦ�P؈q�σkj�3�K�,���"������Sbu��s|MQ�Dd��Xˠ�6��Թ록������0��V�BZp�ma^^jvBC��֍���*���\'4x��B����Y�%\��Z����s�Ah,��˺?��O���?����yȧ�8E�뛀��6#�Q���tb���̊��HG-]��<�)���yM��� ���&NK]��:ǲ��tbm����~���=O��c4� �-/�@XQ	c�,��(�Eě4��\ a�Ze;S ]��h(�$�t��HeeZFz��fE� ���^a�<ͯ˩%jR⽨����6��U�ބN��y�N<�;;M�[��i�н���\��R+5	΁JAA�-[w?�����S�'����yIi��S)^?�Wt�ԧ#?�a<3V�n��E4�S����	Ԡ.������=)q��X�i���v�Cu�A�fJX#i��7V)h�~%d/�F����.�F��(��f"1NI������NlW��x�)=��xM{�LNjAM�+ӯ?rM0�� z��D��J�O���:���IcX����وT|��T��f� �G���ZB5��H��KkCIaF����.��gZ���bH���!-��;.+��3-�Tk�g��L��V���ց$
��t7L�9���줔��x-�[�v�9ӏ�͎��JQ�b��"��(�Mop��⿽���d�z�y03Ռ~�:qc�L��@��]��8%�ǒ4휦w�B��$�k'g��w��W�c�xhҥ~��y��>��J��N�g?�Yd1�V�'��Ԭ��%�T�^�߻�sH�{}���Ru��m^�-�Ȁ�Y\�F�!���3��S?|���s���ֺ#� �P�t��Uj����Jý�;���+�!�x��pN\�dԇ�,V)$Bؖ���}vc/�$�����
�S�&�˯I�#�\�8+�7]��8)n��6J�y�l�,���p�+G�3�xj���F�⑐f�4�dƆ����'�]X����L	܅Xɤ򖪊s�p�CR =�h0�g���L����8���f�7������,��¨��֭�v�~�O���t��ݾ��o�cSc�Fiw��,2�KK������3��'�(���!�\��kE'ZKZ-/�3��$ui�D�3�LJ���Da�.��7y������=�:9|�\������ٔ���\H�)BA)�:l*K"$�5xso�Uyxأ��E4a��Q���4��A	�� ����ܻd>d##�jD�(�)/��q�a*x���TQ�GzUj7�ɒ'�7�
m�o�c��&��L̓P����hSZ9A�)Jt�C#�lnsX9-�>Rt��@���H���F#:+�2PTW�n�{=�w��FϮ���_ժ���v�_�~��֫�ԃp�'z���N2��gt�I����T�e�<T�j[Ϻ�IV(1�q(ؑ4@���S��C�W~�>���GA�oe�>�+)�
$��>e��Fª�F��e�N/+�IbmZ*���O.�����X� �7�����+�x�Ł�kX�be���A�\���?ɹF�t�E��:j������<u7A�G��WB�Nα�~�PB{��hqq�{Z��^�a��R~�k� DV�g��Sv�}�<Tn0�b�b�t���`]��BYw�D�4�H�ɩ����'��Rmܛ��h�y ?�PP^[�eo'��]p�M�e54��k뮫�Sd�F����T����uXIVTQdY�d�
P��h8!��#�7>���]�G�ٽ��G�ϯ���H8O�Z��?���xH3^��2O#~��}�}���:=��ktb�&�~,�2T�"��%6��&*��tڐ<�:�R}���b�
�V.���N�#}����M[����m]�x .�qeݼbKiG���m^][FX����mjp�!��,x�2P*�J�[��T����'nR+\RU�)�rX��3&v�{��62�݇N�.����Op���۪?ۮ�qJ�`�'��H.N��5�Q��P���V~a���Ĳ*�g��e~</뽜�*Z�����g��";QwH�(���M�şƞ�6�����iC�2�$q��@�(�^Zs!��"���p`d�؈j�����N4�uy�,U��ll���ZJ&(�#t+��~��B2����ハ-�Ď�#���ڸ|�\v�Ҥ~��tڨk�B �N��^Y�r2�(i�]Zi�[]R�Fەi{�t�?�������	L2'�7��@Bk.k�F�Eq��kM
��r�NB�v��F�cZ^�"��Җ0�R��i��*�T+�b�e��G=����>��(���+��p �aU�N�B�ti�U B�����F�VlPl�ρfnq;���!�{'�x��
iN|B}�|�H�9d?u=W$�RA�_���:T��;�g]����8vcW��ْLk�ƨ��觮��l�OS�'��~NX���j� ��R�P��,A��_"��1�»Z���Kأ��U�mi��h4��;5)c���4�@]�:}�}�}�V�Q|Ȗ)Ak>�V�P�)e���x�Y�M�N�Y���\�"����[�	a�{�s��Ƥ(+.HH��W���ˈa�v3��D�����My ��3�27_�E[���$p}��I�=((�5 �cP�'I�ٗoN�y���Ԙ�l�x��7У��}z����ӟ��l�E`x�7{�����.��p,{�e?4�T�WA�ðl�~~�:{2��_�G��#4�0�bDJiY� �n@�E���F	�p%'^(��J�Z��R ���.5i�33ņ�S�p�G�`"���:N�T�4��i�롲xv����H�Gq��}�j�Y��K��Z��F&��Yo���7ڀ��4�)*s\�F�=�Xak$������b��%�]4JѹJ�R-�ueV��O�|�̼��ib��7�/�;���v��
��L4,@m���`��w�[5�k�������4gS*�ʥ=IzuV��譍M�&�u@��7[�ȑ'�"�^����F6P��A���H39��>�/MW���H(���{�֮�~R����$G����s�wʿ[�1��Ɲ>&pu���ဿ���B:g=��G�=ȩ/���`G��["pͧ�4�����>�=m(���*��ɉ���?��-{�T%���Ts.���!戥�����P=�"Ч1�Ѫ�b̓�
�Ag@�,��2L�Ӊ��yӂ0~^>]�U�+�`�0{��Ɔ���d��5����ZOh#{�;[�ۧ���g=�n�C{�����;��4�e��H����iff��>�%�7�Z��Ԭ��7�bM8 8viL_Ey=Ӟp����򭇆��<��^a�T
[*4���UIk�!�dfQ�|�p�Z��t�	��pz�V��h}sWZ� Sg$U�MvsN�,�ϲ`�vD�_�E�߻�:��:s|�uĔ��i�z�7��Q �naHv�ӏ�r*H.}g#q�k�p��x��$�k�U�u:�u�KA:��УZɣF�F�'V��+ǎ%��r���vv7i~a�v�u�Z5%�� �2���`��걉������5,�f�X�91"��L���J
���I��z��/3M,R���S62>ʹZ|��I���9<��lwwT	+�P��J��34�z/�,���W��U6
36̞�֌�8��(-,�7Į��Em��g��$��|����o��ߦ�v�o�6V�Y��Z��`� ��a����DZ��85�%+���4�6啦���Bկ+����fdB8l�J��N8�D#�*��:BV'�ej�`le�AB��9z�]b��j�h	�u�H�c>�̫t�l Vץq	)8��LB����?W��+������TV D�L�O��:\���o�[�1�\s������[P��cp��:ͷ�T⹻r�5�k�����Y�������KH�N�jv"����J*uS1��w��S!�8N�'�lP֪o�"TW� �R|Еg�D��_�F+h2Mx��n��ᒀ�""#�?�ND[�	r��a��g���9>�f����s��k��nR=��F �۔=f�BD��*�̖T-~��ͯu����ݼ����K7����)���v>��̺;��^4�?o2�%�Iz)<�נx
�
�Wύ��;�zT4�a�o B�̨�/i�XB��{��>�Dg�B�MHo�g��}Z�w�>�3t����Z�w�&�M����aW�_��㧀S�>A�5O"j�ƫd� �X_��G��F��C����=ׇcr!M��,�p7�&C6�;������Ą���@�a���9O��Zc�]�.-?F�}�#T�M^g#�qЦ~����l=�f��h��k|�ݾ�2=x�q�LE{��KU,�rP��tNK�qQ<D�����P���z��ʘ�ڮ.@�T�V�>e|d3���JU�A�԰��A�<��C-�*>���0�letᔠ�-���NO�i���?GK'/P�y��3�������l/C�ċ�!�� �U��"T��&�&���9�#j�ߢ����ts#���st�=��{_��������5��*P^�y\*�M��Pٸ���n�hP @v^\�1��ϰ*;T���]���G[���H�p.�cO���iHL��#DQ����%40Jz8J�rem��]8ǋѣ/�]Ǆ��W��loXCR�]V!�������k�����&���J�4u���|g}�y��L�d%)d�[7�'߿+)��\�I����"��������+�4�eU��gk]�^��2����,��=�i,��X����Ry��]��O��}Dg�NA2�Q�T�\�HB��HN_��`�R��0�~�����d�!�b�_,��YK�D���%�����VpXI� Ц��q��S��|��f�#ɘőx:-=�6��s��`������:��iVzN`�o)lezR\���4+���0����.U�%z�/Rw��V.����9Z�i��mIĺ	�i? ����a*a�M�� цD��� ���O�O�T�x@��N&�^Uӊ T��	��|��$��@��3��������׿M��i��Y���H��?�B�U��i�G��V�Ш?@���@2 ��K՛6`ޕ�"ܸ[�oW�|s��ۯ�x(?��lZ�X��p@�˴��I_��t��)JO7�Z��%����
x��d��e<y�,u�c�]~���d�	H�F޹��u�9��5�ҝ0.���d�y��Rl��W�Z�}�#@nC�'��%9�ɵ���[��ʴ�4"<�$��y]	��>�^�Ʈ{����q�����x�C�H寮��ٕE޴�H�=��Y��:���J˳��Ez�zD�4TIZ�fvh�Ӡ|�z�ׁ��x٣�'��c�BO��ߢ�����qH�N��cK���7jt8�jP�ݙ�Լ6'��cf3��J�eF�ӵ(�:���ATg����0����֓4����z�]͙,���1�KW�Pu�A�|�*-���iSC�ƃ�.qAH�����!?|�F�V%KMI'�>G�d��$�w��Q�����7���S���G���g(T{���t��5��^�P�Z���k�t}}�x�`	 ��`٧Ź%���N뻷�{�卲�M=!��1�0C��X�j���i'����9HKJ.Ui>$$wR��*��z�<`ݩ�t��dvm��12]����.#Ef%4�V�߉������k���--��`H��z~�k���A��>�2�J�O��v�Q���R�V���&���T#��+��pR"�-Kt��w��)ѵW_��[�i�R��@������ֵ�����=����G���~��F�D'#q�P�\�B}Vw_��ӌ�Ɩ�P,��.�*���xy�Z�u7Β��'ı	��D�^aOԧ��+)�E�*�9J�}D/<�<�"�U$?Χ��� b=vG�huT'�qr���N��BT������h���s''�Z�&��J�����@���L�u�G1���N�k�����ߕc�.ET�TX�>�� R�I�a�H;}�n�8 ��J�mQL��
�mgoce���}��� ��/�x��?�x詒TI�^�Mg/�T��q2Ke:�3�#ϷZ$+�'m~�c��B��k�
G�#�e�a��0�ȍ�
�n1�Uy�I�Pz��oܢ�Wn�ډ���Ga9G�nޠ۷o�&��C�.����g٧zk��G:Z5�w���	��M�S{�YK<�yGϖ@�xI6��f=�.����|�g�Y}�N��(��A�.��,}�+_�'>�qz����4������o�H���n�KU�-�ě���IBCQg��0�4j�w^>f���"kޘ��P㋉K6�o�>�T6M0G4ڶ�/Sѿ4��PgC �j�A�3s|��l��hv~��V�����e��V���^��~4V(�/�|�֎���G�S��{O��d�L~��;�=��ҙ?�,�;���	٦�t��G&XNY\�˳��:���7 
s�O�v��vv�v��|4�n�~���	��{�<ڌW�ӵ���ܮ�s�	V��i��迍@&�11BՊ�2���}N`i�B5�[�ȂJ,�!B���h�c��o��<{C�ϟ���ש}�:�49l��)e��w�C�.��0RjRs�$O]��Z�	|�h�����A��z��BB�pRX����@�� h�8��d�;dC�<N��&=����ƽ�����_�}�;ߦs�z��_�{��?�<���U~��CZ;���8�u�x<�&�r��� +�<X�wե:�DR��TS�5.�����Q��!\(=O��F���X�qBt����̙5Z=�J�\����Yy�|�Fu�5�S�����Q��jO ZQE��	+�Ju��W@�I?�k����Ds��I~�v*z��6���?o����_`��m�`<춎��:�PDuｧi�`�]��Li��n����F�؄B��t���� QqYU�V�K\b ���*q�u2�#js�P�"U�BR���e�;H��X~PX�e�M��F�/�"����]~�
�=� }���.~����3��S|��'NS�=�����1�t������ôv�����Hy��پD�ݗ���vw����E�B�{�v����3�诨j��^���A~��s'��t?o�%j����@T�+^��Vg��������uz�+ר���#�>N�7n�s�~�._�	y�����i6f0�������#dB߼�G�ӡ%�3d�2j�y��9OVd+��J��}l�b)َԳ�!�E�� �K�347� ٥����M{Z�"(	H֚�xu�?�������t��(�c� 
.B'QN/~cWB;�_��{S�4#�y���$��xoC��J\{��֖ٚ� 
�QoB��Z�`.B_�=��0��N�´إV}%TyګS��PQ]��� ~&��"[�'��ĺpu-8lE=����`��MJ��>���7�i��Mm�Ŀ���.���mn�	m���>��r����{��X8˟ݥ���vn>G7�<E3#6�m�V��0ԫh ��XDT��x
_GnU07�č�J�Fl\w;�h��*�̞���"]z�:�ݤ�˫���>A33}�+N���_е���g>�7�����۴��*ݺ�IO|�	�ܻ{{�Y���n�g����1Z�AާZ�jl��W��0�|�d{!ؙ���W����cjV�x�LhP���6�Y�b�ku���v��`U�E1פ�����%�����g^��<0OTA���4������Vwf�1w�2i-�L�����r����"�dJ�Gˈ�&�l�]π���&��6#�73�B�%�����xVʽ���!p�+��J�^�E�=�k|�m首�v'z�g��,_"�D6�$me�N &u�2	V�Y����J-iB�|�P�YK��Z�ݳd!(3��I�k?�|Ȣ�ܰ��X�n�Ћ����>?���w��&�8���i��J�È�z@�V������?JgΞG�KW����[4���B)��η���p�J81�=�<��P�U�%O����������ל_4�wh��<m]nSz����t�}���ߧ�@=���}���F��E���o�g>���?�{?/�������"jD��8D\�Ic��r|?ˮ`]Z�	%Θ�NU:O+�;Ü5q�L` ,0��.(���BQ�0&,� ��?w�66wi0�Bo�̿��d��ZT�� p�B�6R�r���Z�}�y^�mz��G�2�E)�H�����5������d)HY&�QmP�� G�h���v6����gϏ��Z�Ej:���wĨh|��~n�	j}����1�p��"5��Wa�S�4�)U㏲i��w�D�O	x�YKoq�e-�'Sm���!���/�KϾ���~�=}���-�� ����)��>ݸq��NpH̞�O���W����7���Jl٠�4��ޅL��+���}<@�Aкp,>��d��B��3��`��Jͬ5�pР�=����ھN�_�AgN�DF��_��/ߦ�����?�i��O}����3����އ0������P�p�K��o���(��,#���9Ī��=7�P�+4�>� ��B�i,�fe�����t�=��"��6c�q^8"<v�lM����}�߱��ıT�����E:�|s/�8DJ>�B��m�74Gx�O�ŵ=�EL��;�HvZ���{�QHE�.A��ØO��4�OA����,.Е˗i��<�,����,ԫE�cw�MңARλ|
/�jh�W.Y�"�2��81�ޞL�xn��BhE��X��RՖL�l9�>� �,%#5
ri�bB���o��qo@7�� ����hne�vv6��=����Y���d���U9���:v|���/�`�6�����*5BL]O���
ʡ�㑐���%�@xh/���Ddj	oAZP�a:dO�ܚ�Ag���=�F�Ns�R/����u:�p��Ww��>J���O����M~�{���}�q�������A���ɟe��ȝ���Kջ\#$O3�l�aH<c^&�dޭ[-֚V���F:�'{5�l���3.��`��i�?�"�}�l�c�����o�7gvf�٤�g9��ĮW�����p�ц����qg�T��W/)3���=�z��G�I�(X�o�P�6��ʄ�ZᐁOCQ��*��l�hyq�n����b�X�4Et����-`���������Cr�(���⭧i��@I�Y��	��� E�kJ1��Rc�:`Xݵ�Q��O"�חi�v�e^�|�v�w�G?@'zj4���q̱M��o�ѩKT��$�s��^��p�봶�bO��~��V���C��	M����&������.�hlD	9<I�!�� f�������"zy�J��2=��%>(t����D�}����:�Ð���>O����>=���/~���@��.�8��i�T�x�"�:ں©�|�)wu��ߛ����^�<@���)��d����I-%�����/��ߣ��s�����&�����E�s�Nlm��r�*�!~�ΜX�ޕ���hff�6ق�%k�F5~M�\~[�O��d*�W���|F_�~?�%Ȧ��2Eۣ��A�.����b:U�1ѯs��[0&e���G�׻j��7ܵ��)�ԁ���.��RW0���~S�Cywx^8r�z��R��y!���?���\b���]>����m$m�8.76?Rf���!���!�J�0Y�b@b�R���EN��jM�?G�R^�Roۺ O}�U����:mm�у?J�z��H{���J���:}�3�v�_�K/=K��NS4Х�Oᘽ��I�	��#�E�ImJ�Q��6L%�\�l�'�������5�8f�V�#���(ټR �-y�_|�&��ܤ�/^�=�S��?����������O�ax���56����&̭r�FT�5���Q�����I���g��g^�oD/��U�2=P��|��A����E�GT�	���#��IpED�.���sp#�9�Hܦ�KP��%���GC��˖�E���<&�̩S�|�Ff��ȇ;���/�k�W]��6����^���T3�����W�3 ����&����mJJu�x����H\�E��� �"[���s�K^'x���je�8x�����p��z��0(�J��CB�ZϳZy�p5�P���p�<2��i
�*�I��Av�Σ 0鲩��x�kk~u����>^����A�[fx��O��9�#afN�>>1�S��e�u��@A�� �X7%o�V�F��T�����U��h����g_����>I�����K��@O}뛴�~H����K�5ZX��5`/��h,)�4��/s&�������M��Ѵ<����(�8�����VW�D���բ�ڵ��$7�=x�rn]�A�������^�E��&�`�1x������!U�:{�p���/�ڷk�T������[gR9_r���}NB�	���)\���&�G>��U��U��@�(�A� �#����n�}����K���]�*z�6ҀI4и�`D$��}�U�;���B
?Ѳd	ǜ���-�@��\��k�+�Od��wib#���}m.q|��tis�6�w�	^7}:���c*�"����ۡ2��`ء�������F�����d�Պ�����'�#�Mz�j�b5$m	b��uz=j�T(=9O'�����.}�J���_���+���m�~�)��_|�A�^~�eJ�?N�Ǘin�a]�C8޾e4hZ��G�|�������ԵM)}�C����V`ɖ�̥���`q���n��|�ʫ<a� �IN���� Jۨ��ȶ8vBN��˯_�ǟ8�x��7��w�r��;_9�ǌd]������J��!�h)�:{��̬d�D�~�'I�mooKJ
)3߄G+�O�>�*l���B��1{zR�T��ҫƨK�Ŷ�#۴�Mr��s��x���}�������Z)j.^C@)�&>�Kx�Д��}���ݽ���:v��������v�.��
��2�����i��bЂBh�����砼:1!��cTB��!5�Jt��)��v{���s_�O}�����n?���D���'���/�#m�o���&5�O�p�.l-�};�bXkV`L:ޞU��6ޙ�i��Ɂ�^�[�Ә[s�ą���L0I[[]�J��GAR��z�Amv�$�w���$bk�R��[�:��*e��5u]��7��9Oq�'zy��@ߨ�g����;����yǦ���0źt,LW:{�<�#wbM{*G؜))��l�0��X��}Z[��vw���^h��[�;�=��{��xI�Q�GU3@l�Y/�����s��6�<�t�.��@hi��"]�=J'�o�K�/�g"AYvϒ$��]y�Y��F|/[;�������Ю�A�Na�0�M7jӀ_{�՗!�;7��%aRPR6�zܪI��ܚhZ��<����X�͋��DN�ߓ�|�#�Yd�U��1�9W��NP�=�^x�7����]�������瞥���~�����K�r�-���7�_��K299&G
�#��q���XY��A�6ͽ�_`52N<�:i�$�
[���}b;@.�g��K���^�ۈEP����+(]�+4���VC��w�^�(N�C^��-JE�l��d½�}�h�ߩ+��������7;��R���~��b�	8B���=�۷��Nr�R+��˷�c��Ͳ� �\�Ȇiw�0T��Wȯ���(�"36��$C��s)��R�Ta�*�M֟�ԫ�-����[�Wql&�K�(�ڮH��:b�w��{�����B:���XD��^���]:��jԫ8=���pVX���v�v�a2`�p��Z>�1��0�&S�2����:LP�qzn�^��:�6*��/�>������U
n�ӿ��ߠ����t���u�
�:����4���v���IsFr1]�[��+O����ܥ��T������D����1��jL?F�ǩ�Mkmm�.^z��ƑSQ� c�=������"�,4h~����]�EN��
n(P�ɍ�V���ِr����)F�{M/�<+b&S�����.գw����̀��M�bd��
���f���]m�7�z����c�LRDwlm�C��qJ	�#��Z��=��wC�mq���)b��۱np�H���@]�V�b�^�ƄNԮͼ_H�Y*����C�}s�8?�v��vpg��8�o5��4�>���{l��,M�#�h�%#���@��8:}S��]�!�.��k%Wt�jh��e���9��QҦw?t���:��ڥ���A�ٯ���~���CO~�t�����mL
�ͫ�FE&-I�>0u�BrT/*Q���p9�Uq=�c+�l�6U�t�����)jQ��+Րj~H��1;G7o��h���MT��}i��VH�b$�2�0ͪ�#�[q) D�ÊPÅ!V��.��!7sN�-<��2�p���u9�Y��1y��H�v;CZ�[��O�<�^���N��+ �:�.�/.S���F7Ǐ���Q
>K�٘
{tNĥO@�uq��#����D���a�if���ޚd��(��`B]Eb��>��/�G7�]d_���P���������/��{O���L��T����#^GC�vX�����?�>(4Mb%}ρ��4��E�ml4��[c��yTk�(\e4惴J�O���A�.�ށ����?C��?��h�����������9ޏ���1��[챥6�j�'��8��`���6?���H_{N���.+fk�?UA=�D�_�ȲS���W(.y�����@��]�/�E�ql®��pQ���!%��6�_��'��TM���r9��n��O���/�I8H�%��:�\f1�]���ӄĺ�9ݱ���-�ܾi��K�&o���}��.Ď�T~�,�6�0u�j�?ee�T2b����f���L{{�tlu��W�Sm�8�*�?GWv��c>�w�v��xՋ�{�����7/��R��S�� �m�T�/u��ŋ�:40t\�A)�R��i8��N�Ї f���i��C�k�4ߨQ��R�%�r��9{�ac�"�hI��H��;�g�M����Htٰ,��yv�����q1�3���jau�:i�Q�p���< �x���g���*�8�{���9�G��?��>�U:��������I��{��:�mZ[^���!�/-����M�<�ՠ�sA�kGgx��\Rwi�h�ULch��e�Xaj���M	��lӃ�@�㮝8�q@C�dss5���]T��*e#���\�3�K������2a�Ϯ�в�h�&a��U���'�N�[ё�[����G6�e3�����Β� ����;BY�%)��I\]bϠ���%�)��,�a_;��:��X/�q�R���9�߿�F�8ö�<�F=h��t! 4Z[=�Z��FZ�%�4�����h̩K���Y�A��������T0�ا����/=�}��l�>���.o�KV
���`����;D� }e��hH!]�a'_(̛�5xZ�a��<��ȗ*� ﵩB��KmN�A�^��u��[�e%U���R���ڣ�/^Cs\i�������|% %`�����G��+O�����=Q�f��Ve�R��&�4���H���g�ǐz�y]�A=��U�2:1;��iSٻ<�B��ud�q�r-�`{k�O�>&�V�a���Hjm� ��:��x�Z�Yv�"��bx�ƫ��9��w����^wC��)Cq�:��M#�7 '���{/;��@%?����V�{jҜ
nz�I�Z��P��@JS2Q|lI��!�AE�0˖��j�������}��A�=|�2E%��f-0�����N7���s`�{�m$��ܳ��W�^�8q���8�aH�p����L�!H<���K(+*���������k[g�I2�0���Ne��;O��4�n؞}vj\G�"��U�9t����Q���uo�S�_���fC���Q9���7��s��7�A������)̌��_d9�ݲ>�z������Ş�"-�F84Ξ���찆9ފtn�J꜋%��6Ǯ��;G�o|�O#�F�N��?{�dI�]�]_�:"eeV�ʪ���B�!�H���bI�����Ѹ�ΎF4,hr�� ����jQ]Ze��p�{ν���Ȭ���o$*3��w����wŹ眜j,33/�����2<�pW��͙P`IK�r�L]���~���K_���O=������|���x���jCV<x�ã}y�y��d�։h]�%���=��/�!���}���1W} k���r{���'"&R�|c��x�z(��y�����L�q�����,�e4���(�����z��lɣѩn8벫aҤP�W=�����p /ݽ+q#&j�\Z�a$q�n���EU5+��cl?7ȿ_��(q㳈<^�g
�K����#��H�r��颠a���=�u��|��C����[��Fg2���gY��\��I_Zۧ�w�*q.�3�_�{�����j,�H�2Z�d��������*���Lq�~��hm�}�6���}����~������5e���������E�MI�\��Gj	�l�ڒI��	0Зm}�L�2�����S��'/��	�'�H�A��|��ڣx��%U�p� ���ᓬ~���?�.��ʳ_���ϙZb���p��s�Q��ÍV��� cFV�V'���k��n24
Ղ�+�$�J��L��Y�+�*����;����]jxR��K]��2�&�-�g��%��lJ��T(c��n��f��X���=2P�4Tj�zr���m�#Zc��STG��2�o�Ԋ���8�Pȅ,�bT���HDR	��ЪUENL�&����Ñ�N߆�SoT�{X��+ ΅p�μ^��d08�O?�\���[� [ ���7wek�'���}�'���z�kRK�*2I��u���B�V%Y�!DP��@`d��6���@X��y�� �֭/r<�ʎZfp	"F�tGc�2j͘	!Z2�P@s��^���k��/w*{��z }=�� XJ'
:�����	�\G�	q�3��?����#y�!	��4ı��Xl���_�c�o�,�j9P�&���Cٽ�Z���Jdߣ�}R�a�)L��	��FV�� b��G��7$ꍬ�#(E6gS��uQ���j�xt"'���X��	�2r(PԞ���]ߠ�A��}�p/����|Y�$5U��|Yj��\�S�_|��rn��2̥S,ևQx"VJ�L�D�C+Z�������OC�\�d�����=�'��IF��b(��4�ܐ�?�����A���YCVE���	J�� `U�C)��%>�F�E���yE�Gb�i0Ǟ&Y���N5��t��{K-� @�hv��Zi�pG���z]��M�����R��[&H�����+D�_q<-�P�Ӑ$�9c�^B\xb��>�l9����/�4$� ���x\��l
2k��;~�#��#f�Lj�D�������:��u�;?|�������S2+1{�՛�'h@"�����ҋ���aH^\^��Px��J�̭<�<�/X� ��s=�@�S���J�vmTg��	"m2V�c��l*�Re	Pk>̬����w�0N^4����?#d�C�V/B��oL�'{NKή�+���$QE��8���YݹHMӴ�(�c���2>~�f��zJi�����6d�㙜��~e����C&T� O�-ƨ4I������r���J	@2�{��'��,��(	+��&�O��d�	x5X�����mI����쌓���J/4�ftoG�X�ق]o�zG������Nw�m�)G={�t��g�<�D�f�_�z�$�ҏ �Zr�np�j��Ƭc��r>�|��������(����=f��� �� f�(�����wYF��1I��j��%1�kZ'�rH,�tM)p�q+^�d�����"��q>����������������~�JN@��ٙi��'� ��z��]�zn����w�t�0��q!�>��'�ٖ"�!Ѻ|�Q����φ�b�<:\P?2���l6��"��okX���Y]����ߐ��P��QM�"�\9Ǚ�$�<��oh(
{�(��=����%���1�Og�Q�����E��O�I���mu���p�G�Zss�ͽ���tf��Ṍ�w�MC�l{�*�\J�����V�LGID* ,�@
],���r��dI�Ldy�r%û2x�P��9+9�P^Y�:�|mHZU�ƫ������ǅ��y�{�-]e�����e�_>%[28)��b��&i�x�R���j�����k�Ѱ�Rih�~>�T��A(ħ�M",�
q���N7=2/"�fy읶���|N����|���;1�a ;wGg<�	Th���x�V��Ɓ��Wo^�2@
%��DR���/X.�.(�-n�<"�u�����q9B���]���Z�\a��{(���.�w�u�>��;�PIA�AО�j9D��d���e�����i���k��P������G�7^�zB�#v8;����f���X�e���Ͻ����N�\K��u�*�S/���׮nw�*��[��MRc����/���[k�� iM��jI��nw��	��n(��Hh��x�P\����]��	P�џ`pė�{��<-��Ly5qG�{G]PǩqR�+EaQ�� 5����\�>���xE>;�q7��4+,.EE�S�6���^�t*��ʺ�Q�(�BVg�D�/�gD ��X�J�u�@��1�Ld�&25`[�;�*��Lt�!4"Z�z�䡕x���<��"E�@�gd�*/�?���'Y-����Y��A���N*�%g�]>no�1ƹ�Lᐛ,SC��hWC����SuÉ��}'
�3�����:���K,+-��.��@mƲ�Z�����m����X9/�Եش`�z���%�h *c��с|'��~x�[ݎ�@5
�^���^����w��u)f�6�����4�ԟ���y	[��Uv�R�
�p)x��y�{.�%{_I����܇�զy�~qO��t2��\c��rD�a2^�6f6��Bӄ����އw协��C܇dWr)��R��U��ͫ��yU�(�\�7��5{>��]���W$e�3���eYU������P�N��( ���/�7$��X�TJ$����ޚ�	�@$R�v�Vݾˍ-�rR��`���&�khQ�_��Bl�z��VWÿ{F�� �yڨ�-����Hڤi,h(����"Zݤ�9Yz��'�+��!��e��r8C�z�T8���M���ʋ��K/��#+?��;@S�zs�[��H���K�r�՗d8�s�1�J�K�ȅ�?q=�@<�v�8Ԩ�c}��{W�^q�7�'��S��,�E��m�_c��p�c���F$�Ib�q��\n�sc?�;���)�k����J�tf��~0�
�VtIi���)�T��y
)�K&Fѭ���}0)�\���d`Y�T��΁YX5��ڰ�ba4Ԙ�<�{2�ڞ�;��g~6�]�*aK�l9V�S�_�\-~rID�:"��K��8��6nElJrƏTr!�ׄl�&O�OGP��P��*d��Xo�n]��L��ȿ��{�o����[�l%T��nX�D���(^y�%��d����y��ó@��_��
	o��R���KV���b�d,z��K��G��pt&�NM�QTK]��Ҡ��e�<���毽N�3�3*T��_��<�U��َ����;~@�+�m��'�#�xB/�c����?���Y�>�F�<����`;N��8DoW�<��-0���y,��P!���Tk30M�[^�Ʋ�ѕvW_��HNO�u1Τ����&���jk��G�p�I	_v�/"^>����57�C��02��_��H^)(���5�@���j��i�|���rrzD(*0`��P0��[!^Ꙭ� ^~����Y
���a�33yhQ����:Q#�=��(C���cCQT^^AÁ{�I^jz��є$8���''��fIѩ�����E1eٖp����B��ta����ҽ�L�3���`��\z<���埨��7�%�&
v��DD/��^�򋂚���L>}����ޑ��="�j�Řkkrr��7�qdZ���-QC���r6�L��Z̰���Hl4�g=.��7�e���+?��>��'�x����p�e��Uy���؀����.�޼t2���܍*@�^�+�9@R9�wR�10ib�� 6����IUx���Ȍ\ ��$�0e.hMp�#U���2��Z.��k�U��>B�"j���zB�a����kk�������l��s�<	(g�� �p�`5J��\�2�E�v��T^������ƒ��t.N{���c�B����F��iͪLw�U}1�C�kQv:zn]�޸N X�׳�p��WD��es�K����})bIM��h{�O�[�|$�1��,�DL��V ��\�'[��y�����H�Z�M����w�4s&`��M��G77�[w��	wȄ�x~�xt���7O�<v���[����V2~��(�"�����pޓ�N�6�US����}�=K����,=9r�����I"��'u���ͥ�6'`�0",�a`�Pi
��"spQa<��,[R?��Z���3�} �K�U���]m�A�����Sf��e���Q�c��H<[�bB���t6R�xu�!yc	}+w?�����ൌd7�.^�
��J��.]{<CP�L z_�cF������e��I��S�:�QS�6i{Ґr4���IhBU��V�cD��n��UW�O�"Q,���d�"BΤ��a-�}�r�����&LѬ�&��l�n~<| ݭ�+���G"��hqRN��t�kj	���O'|xĳ�A�:��r3��K2�f��>}��ǯv�o����j�o��)�.s��d�ʦ>�Q�d",��c�1�Nu~6�Fғ�x�
J���_S�?<�2�}H<�9�*��3[\��aIm�%�9
e�E���G�|b����$+2o���N�G�CzY�_��0aUlܷ�($/���2�A&�,.x�]�a��3I�� �ase��Qy!�%���s,e�
�N�{,8/�6yxӬ  �{��y#e:�Xlj��P��|��9p'�E�֮X?��7Tط��HIu]��,9b�4�l��Ī��'70C�	W��˷Ů[$�X�/�p/D�^���ѡ\;;����������_�� 'Q�#���贛K�qR��΋f��i6�F6��n��ib1*DR��^�|�����=�R�a�$�����U#Vj�_w�WW��uT�;�֘�6�>Q8.�2�x�P<�zĲLP{VB��.��.2�� yX2C�����s�Ll��]l:ɼ�K_�aVN�>��I Ԟ�e.�`܎��\I	��7�P�k�g������ySW�b9�|�ax�e�^$�JRP_k����d,�.����,�.��:-�e�j�X�w$�/��f��Ľ "��k�G��O��R�1�eN�E���x�R���s��&YP�f��z� ~fէL��M�Y�;�ή% H�4(?�q�u�֯G�\�"�|"��ꍟ=x$�<���!(�m�B�^�V=�牼�Yr���Jn$��{�T%oK�
�;���3IAľ�lDx��o��L� q��	T^�uۡ���������X�mQ��d��Z̬��sT=��ߏ���2������>B��,��	-��9�~��pp�O�$�	]w�ăɚ��X���N��Dx� ��:2��*��QCϒ��CH����Bg�ܬǬ|�3�:����J���S�0Q�|�'=��K���B��3}�͉;�#c�%)��3T7*e}g��,����yB�n:��+]�^��Ʌ�pJ�R��1��w��a%���֝��������|dmVK:�JO	����MW�NWl�[��e2:'��"SC�,e
�hW����U)��-L������U;��u��KXz�z5�Bb�n8X��㓩�@[����T�'ǎ��OMs�����B���ov�dc}]x�;؄��	�@r3��r�\�j�c���ŵh�o��o�H<ӱj"o;~�}�|<���cf��粻ݖk{:�"	r�]�ȷ��;\q@�QM��A�tl�+'�z�HF��Wu���d*:˨�M(2�3��re0�Fvj��y:f��sJ�O|� J�Փh�*��Q/"wpP}tA����nZ�����^����>��t���r�`r�½����e<rf�l�Y�*�X�Y�2�$a.�V��A�y���rBX���Ò�b>g'��ږ�?8���ޫ�m�����z}�v4�L��ݧ��:�T��E镰,X+��翼�ġr�м��4�OKL�Q]������SX�H�Q���q�͛�|��'r�H�'��Ha	��묱���uQK����=N��\�[���b�p���k'��_e���g��y���*�ԣ,�v���I5f}x��T(����u'�?�K{{�d!B; �j��s*�䅛w䧟|��n����x&�����zm���Km9�����p�%N+V��Z��d��g��k��!I���B]o�PЛа��P3��qiC�Э�5����!_C'/���}�R� ����
�g��#[�Vn�]�v	4��lK� O�U�j�Y��hP�c��8�L-�t^�A@o
*��Ar�Id��D�F����ɝ7��}��g�����[�������N"�f����֝=�2�_:����V�|U��bO��OQ�ރ���E��0y���	WG���cT$��o�-/�pC��99 ؂J�	"'#�⮭��	�|�h��HVr'
�8˴��.��"��*
OܕW�������O���Si�:�/�`�p�޻��\X����]U�V���3b�:�(�/�j�MX��5hv-I���lD���#g4�tދ��M�ˡ��dL�(LRx~P��l�%t���5s!���ēoXx�?ZT����(<��z����n��w6�u{�=�C���Dڭ.ÊV��{udMC؃#�h�1]wVO"��V�O��A0n�W$ h26/���Ą�
k�>[th�"Ұ,ي��Jʶ�y/��2�, O�Y���pp#zI�����RC˶��/���!��!�e<�o���^�u�!5?RP,�Ҵ��
|xt`|�JSKϽJQ:�I
qN�\�cx����eH��WŒ3���3$X�?0�l%���m���jݎ�asoL%9I��Z�1�"uW���eskS��\]�3�ɳ��`BF��8�Qy�PUqaxĀ�y��i�$��$�ȭ_�|tUj���ܱ��ꚞ��"�k�n���V˸��O���XNNL�a�;M&�RN\o�k�r�|�>���&%]�Unf��*b��n�{�sls|"k�5�N���D�X���|�����1y3z���ȣ�"z�j�G�4FL�ZC��=���3���%��\1�^⫹.g��#��H,���˼ڱ?GX���w 1?ӿ#�CF��j�3�����+_��Ͽyg�i�±�ٕ��s9;;b�ĪB�J�E&V�[�G�\�póX�=+��ix��)SmV1�%�Ŕ_~�@ݠ-y���W_�/>�1�l��8���`ANcr�I[���*\����R��TcV^��X���$~�g0
��˪ �W���ِ�K'}�����$2^L4n���TP�F=Y��uJd�2{��oo]�	��n*T�����[��{�f\��`읍D��U:e�LM��GU5�PR+��sP.`9B�I�s$7�oj~�u9�?�����Z7w֥��Ǥ^�ӑ/�ș�OG��F%նx�$ ��#�8ʑ���AD<'1X����2{��<�P<�EfJ��LJǤXX�12���]k�4��YV�!<�ܡz@�󉆈gr��7���������ֺפ�nȻ��|ĕk=�u�5&6�9Q�-̗�n��U��*\'VhJo�����9""��6��3��Z��f{�_ʣө���ܢ^bZ��rL�o�S��ڀae���r{���h���z��L����!?�F��we4.�9���.�����_ݗw��zo�jJ�,�k-�������%�Ƴ1:���˘d�Jjlُ�����-�Z8o@a��z�_6�+�.Nɵ����5|���2[Wn��Gd���si*�h]�]Y��=�-�������F��:@��e^�A��h���pY�J���d�4�NU�BR�Ո �c+oFƸ�D���.�ب�1X���ǟ���@�����Sc>?��L�Q�?��>	�76:R�IT��ؽ�Ҥ�H��wQ����a�!a<���꽆Ĳ��c!�tiO�����_�uGY�g_�ސ��u��}_�� ��T��5�7,ƪ�0b�%5p�߉R��!S}�h&Z�N��򪑈�������^|+X�'_���,�W&C/�I�ʧW3��λ|,��C\�a�$KJ"��J�F���F���Y�5��u��;Zj���:_X;B�MM�D��_�ɟ����FJI���=.����uî�Y���_�	X�ش��5�Ed�J@�����_���"Ü��H67�dr>�|v����w�+Ig��4􈥓%$aY�?�����]���bk67�@@kry�QJ!�.�݆�P��0�N6�r��ͰJ�_���@Y�>�7���G�2����H���E:�i�-]Gc9��H�>�LC��^���'�χ2�����-����K~�;�x����m`<r@h`�6EɅ�ns8$�<�����k0l��YS~V�T�t1ǀ�$��h	-p����!���'��p��.H��1$�䩷̍�K;����t��L�0�g �`Y.��rņw��5,~�Gq鿿�#�b\���>�) ��*4��D�BZ�ԸG�'��������lhBI�0U�?�ˣ�盜�.�+nC$�x���'�®;pI�\��YNO�b�ջ��T�|!w�^�������Җ�F,�����y�M���Bf�T� 786�H�V���^P@h��:Q\3Y�G�!u���(L�XX�~��%#�����/Ίhƒg��c�ѕX���N��s��t��t8���s����W�p�>}@�Z����͗�o��L8om@��Rϑu]ͫL���w�>&��}C-��͇��zg3��^F"E��|1� �ۮ_�cf�x&Cu�'�� C�|���TP�K��~�����J��F!]��&�Z�8/�Xp,�?�����X��^���y����8�և2����d[bZ �A� ?���MUÿP��n�:����}Nz�*:y��뭴4%������%Y�C�Ӻ���v]�0���
���|=')�S*�w��#j��}�;2~�@�[=٫���X�yWJ��N�H
u͇ɜ��\�1vڄ��BJGP-;��0J�oH��#IlO&#P�dB*'��:x=���fhHӗ��z����!?�	J�#y��my���rz���3m�R��J{�����󟑺�ʵ=����ˈ+*饓A*N�*����2����%�	 ��=E+�|#����BQ��$Ÿ����J�:Ұa-�΋/��0������$+! g<��صn���5�K�S��7�؍}��/M��x���(��y�w	��ui�rv6e7�֕]�q� \�r$Ssn�����J����)�
�i��֪��D�s�WG8
F�_:�l�b�6��䬯�U��^�+�_J �Cu���v�e�1���3�k�QJ0}�>��2���N��i�M!o����:S��Y���ʰ\��UyR!�
rL0�iJP��F3�y�sV�RǠ S. �=�'��oK���Y���c5��;�Ml��}!~����[�JSC�(�M!���]��;6��We�.���]>�Жo'���m1��V@X������lB���"�n\��+o��޻?���O�����x���7<`-����嗯�T�k40�lj ��3)<�U���Zy���ڧ ���ox��i��磠p�z������7��O�I0L�Y_�K�#�
ڂ��۝��Z�n<*L�Z��&>�h̋��4�z&-Z���c'c1c���FO�$H�xa!�B�"�~鸑h�S![z����E�;z, �Pd�� �	���3��Z���L`��z�>cw�e��P��7�ƭ��їS�$����/�w������f������H�ː�H�{��T��I;Wo�q�S�=�R�crod���87{���ɻ?���}�-��Pi���v&r��d�Y��{�����A�2޸}�Pzr���	+�A�Ҕ�|�+���w�(��!<�j�J؉T<�p��8v54�̐��?8Ә�'[[rt<�>x��7+ə �!)�X������2�.ʡI�0��,_R-V�hULn7��n�~ڱ�3��HT#d��I�Z�,gbi�zSÉ͍�N���O卻o8��y4Iݾv۽�Q���̩�S"2ɤL�2�i��]����R�Jp&�߲7�] ���=>��)�D�������]}�H66�dq:�9��	`#�1�oJ��G��||�ބѵӥg��bҎ���.2��Z%p��%�����,�O�J�B3� r���U�~Eb' � �r�\+ǇGrr|*W�^��:�K�Ѿ���m�Ү����_���?��o��{j�L,��`��"�ZIC�9خ`ْ�A�)|s�ꅩ�Gl�҆hTt�d ���^��N�-�Y��W�O�xO���ѱ|�08)ʙx�Y ��h�����5.��ֵIk�y�L�JVh�V�1�����Zc��������~&�F��8����#(5C`E�DsP���z
�!u�[)�� :/#�
 �RK��M�̢c1xHIbG��.�RrR��<�B�n�s>W���h	����P���L�굂��D=�����d��n�ՙ��øٕ9�& T�|SǢ)��Q�Ϥ?�K�ֺ@'��1���Ĩ��XV
<s/�0U�@�ܰ�c:����<��&Fly�Ġ�R�M�r8�ȧ�W/�&��}U�[,?}�'�B� 9�^Gn�ݑ����o�֍y�ۯ��n��Mx�T�f�w�Μ^qf&0jP9�s/O_��,=��9�U.�i��X
er�XvJ��p���yr�������믾&?���b�Ya�ۖ�Oj�d�X�e��@",!*,A�w�(�a���=����'��_��؄�،j�ڧ�Bnv��ڹ�n�#;[m���\ݑZ�.���j�[�<,y�O�ִ,yl�3�U�c���9@荴F�ܤ��m݅�W������6�:)P��1Lt>�m��Nt.Ӆ�H�-�&��ht"�,A�<I��ɨ?�"�Is㦴�o�X�(��������+"�L��,���V�����H��x�z͐��k�����s*Yn��gA�Z�懼�e��j�|��C�S F�2���}k]�w��ې;7ߐ?��?�3���z�E��Y�q6�Ѫ��Ji���q'��l��Q渺W�<��D�y�[)�\	����9�ȹ)���a	�;u1����J���hoD�U�����O>�*1q�½����X�R�I�[h�ؗ�+{�q�:�M:��G��0腭������n�-U��e��ޓC��C���B3��a���/�������C.�X��7���.��嬽�t17r9R^BfV�u���"U�xJ��,"u�յ�����z{��><�G��-��Z�{�<�ʞ���O�Tc3i2y�Ԍ��z&��4qi��B�n�;�)��\@`�r�N�8�.n��H�aZ��-�6c�ٻy[>�חk7�'��-��BF��K���d��î��\�(:���\�_��g(���2}�@�.�z�c*�؍��1n%H�O
�>�,�����@d��h1`Ccd����m�fO¶���wO'�Os�p$��c�������@���̵���٣pο����\��ʷ�y���v��
;����l��5f(Q��xk��nކpsk�1:~�����r�8��8����zt�/���XZ����������q�K��*��g�����M�#Q���Rwn(�|,��\�v��dX�k ��|�c=���T��O�R�a��Q5o]�����<���c�}	�t9�yV}��;[��R`�k�;��4�k�{��fC���ρ@�f'h�p �� 
��U��d/!_�kp���ἅ3���J��5�Ɵ��6�����9b�;��:�b� �ڭm��O�V&镗���כ��G0ғ��2�k��E�笽"�/L~����X`r��&"ރ�:F��-r��`�,�rU�HPdP�K�z/�%%`�Ѝ�ܟ�H=}�óƆ9Ս~8�ũk������ߕ�^]~���Ui��!,<�����-���0��d�.������&�/��q�1~y�dF�[�Q`e^��f��Br�_�:��~Y676drx"{{{r�ӏ�x�{E�	Yq F�\ߔ�nS�<a)h����X]��`��ϳ,T~&�� �.W3��j�]�_Rv�嬳����R#x�-
98y$;;[�	���[�y!똠��e�v��j�lj�'e+")P������%�Zc9őŵ�eZz�F�f�FHb�a���1V��������._~2���K������Od�=��ݳ0��E��r�;��ؔ��}����Ϗ$�K�\�q��'�Sjz��&.%gΉ����z⑊c�﬉߆�:+͞B{$i˗�>�p}ʍ��m�zx��ϝ�5��k��|�ӿ����仿vW��pS��ߡ�ı�_]�e�����A�K�W�1.�ǘ��$'��Jfy�Ũ6o[$�Soa�D�H�U"h췷�y��b.Ñ�8�1:9"f�����]�Lݧ�M6����:�����B\6�`���Z�8����4�=K��-a~��p�O4��Qݨ6 ��nm����C���˒�:���E���\�3#��#�z�`��QX����Z�$U�VF�-�/3.-�Y5�1'��Le�\����˧?�#��"q����9`&��p�-���ݴ%n�*��j�x��L>�K�|!�w@��Q�c�~>E-"�rz�8��C�Im#���/�:����*C�92h�Á��ȤN�:@�P/����|��F��׍��[�O>�@�y��|��I(�Ee��3��ZjW��A�S���e����, �B_k��R*���}a�-��'ֵ�q�!l!��-������~�=�Ͽ�Bnܸ#��H�$bĔ�4��'C�hL�җ���2��x*c<�Gp{�������x���<��!| �+����B��}����=�����G���)/�x��(�t'''j(�$���шd�̑�%��w~����p�����2���.$.M wj�o�g-��^�:�.�d2�'�.���L�U/�,݉��aB�Rs�
8
粮�t|j�ٓ����-k���.�=u<{�u�;
7����S��:��פ}�������ߊ>�b�@��!٦�������S`(��j`4Ċ�Dt�Q�Ul�$k�vhDCP^a��yAھ��������0��&ۛ��u�dO�<����L?Ӓ�pB�	Fj<�w��my�-J�ej�@S���4Nl��TV;?�̓Ĥ� ʸ�!�;9T݃�I�p�]�Iu�5��Sh���ƈE��b^�xhM-��m5 �v���-+�')��rKYS�\Ͷ�lo�CM$^��K_���[衞�Xl�KF`�};�e�� u�A��[���':1rscK'�H��F{W�U�7�歛���.V��l���ҧ����Gk�	ݼ8 �2�\��h�J������Y�шL�;f�B�7�I��
p	V��;�-�"c?��/�NzG�W���^m�w�>���\�ʚ�G���&������'�Tw�G?�����tt�޲����HR���9+-544�w�H3d�=|��;ҍ�Q�� U�G�8�FOZ�z����on���gr�?��&��:���S,��W^�W_Y�b�Ƥ%��I�Dl�a"��ߥ�1��X�]����̋�(Sd�8!1�A�b_��\
 ����5��dK'�*�rWo��ܗo�/��N�i�z��,ғ'��9))�������"��k�v���\D(^X>�c����_�ģ�c���#�Zg����}�����P'��|��z2�I�l5�0�{���J	m6�37��؋6�8O�
��]��a��mQ�rߍ��άH��K�9�"��[�B���%:l}����˛l7�E%��ГQȩ��>�����諫��Fץ�\������-��a���{j�vNltЌMk��k��ԗ܉����^C����Y[N韏YS5�5DY�L��P���X����!J�X;�A_Ë���5y���'kj+�D�2;����ԕ)���r(k_/���i�  �A	j���8��Vq�F�㺹�gg����D���� �$�s�'ܸvC�?1���ӕ�4� 7v4Vd�0,�P���tzV.�X��,k������,=�h�@y�52߿P�D����F�������CL���MW]��N�r��� >�;2�ݭ^S�b4�N=���1��H oA.���x ���G�-�!@�*`Bp ��aD�w���Z��=͠�T��G<����^-ӱ�`8��u99:e�	��sE�}.��L>���养zO�z_=A��\6���O]�Z&3u�);�F���կ��ԔNcM^���Iv��|�������D,fz������������D��dhqzv&Wwwd��loAA��c[����/��/�Cџ��#ٻzMN54�f��[w��&k����g�'����c��J��q`��X�p��OXK�-�`&�>^�nF�|5�_�2.��r�:e�A�sǩ����If�2�_|��$Yۓ�7��{���~W~���HQk��1��d��J9�S�I�ӑV��߯�Y�Z��zG|�劊.�@�
N��Z>�ŗ�T��Q<���݋�t�DKV�'ރ�T�^U�ߗ/���̅�\�a�E�<�G��iFBd�@�fC>����6Uu�mG�h�#�\�e��S#ޗy��Mc2���O¤��X�}���ei����0b�����]���9�?�����U�`(�
*�|����`p^�|j85�᩼�7����ߐ�+�������E��@w�#��D���Y�R�4��� �\Sc�;�|*����F�����z�y��L>�Pv{-ٿ��]�5: re�}lQb6�ؚ��L�y��be$'j���hp*s]cw�u���m�n�d���6Y�Ъ���5����@Wc�$��ZUz�G61�4���s�p^�bJ�+�`�A�G ����t1���%�k����>Ӹ��lc��7��E�s����-J�A���8k��M���f�&y -]�`.T�2��.mV��b�����{t������c�o� ���:!Kd��ȉ����ɴHw!�V5j���Av���-i�u�M���>�RS쪓�aQ�$Ywt�H`52\�!K���й��ZX��MR�D��@�[=	�?K�t}-���\��A�;f�e�ɪ����'�;o,;׿#i{G�	��e�)�њ��Bg^��P�xr:Q/�G��B7���z5���c�۲�����H�h\��b����&�Fc�Ή�������`���z2�����>�z勁�4�i��rmoO���۲�r��Q!��Y�݋���
J]�]�ƁE_aC3�W��W@�[U+�,)Y��1<��-�D6r�3 F:�K�A���c��rW�vS��]����_���؅t�;k�'��1�JWݶm�Ӊ�����L��`Ս?+�zE��\�1�q�ӎ���=p��2�@�H`����VW�"�L0��z9���_��h�']Ʈ+�����$!���@��6ۼa:���JC.i�]�x+JV���ڨm���_�t�l�J���S�$��#I��&Hn���3���?W��r��oKw�5�vu�^WCu�WrR`(L�2/4�B�a��E|&��C�O�5|��!�J��MR�gǒ}YL�Hr��	��-}Ɠ����ō��|V����k�Ĕ�Є.��������)9.����r��Uubi ��6����Oj�Y���.�Wpizh�r2]��x�9��eY�Ʈ�G��-_����^��dlm�X�9)�m2!�8f���o~�CJ��o����ٕ��ѹBN�*�ɰ/�ф: m(�W�m҈�j�Vu<ɋ�;8B���_i~	�C8�E�Gw9q�s�0�$x�[�C�s���J�Ĩ����ӵ;uk��	��1d��.@^��<�j���Xw �~a ���Mի�I�����J"�<
�D��x8�LG����� צ�p�|�2@�K�jr~��|6�ɵ���o���X>m5!`4j@DFhlBȤϷy�'�١nl�����_h�,�L29=�\��Ո39��R��}�J�g��H�S�a2�}M4,��O�a��l~���)n���[��-���%��P���ĹZ/-߀�|�!;+å������3�Z��W�|E���F��\"A}��ʵ4�s�A���Q��ZK��xQ���_��7�{���g��!�_~.��r �L4>a��j��tջhCBlCNO1,!�1�&v��"
"Qe�'Z��x�W]��0�~�E�,�̋���ǌĪ����+���=�~���Ѐ/ֲ��X::0�}n��j����o��!�ɋ�`�����|#5�Ƌ�x���e5L����rK�a�^kyM���xx�C�7s"qJ *q�1+,Ё@^��Yn��oeҟ�Q#�Q����}# '��|p:���o�˿���K8�jV�9��!��v�28�/��}Y��}����gihx�fr>Nm]k����ښ��;Ͷ�}i��H'��	ᨅ�����C988Q#r��uy�[����&������Ff�p�:,\Hk�����U�x-�~8N��;Bߒx>º��Z�22��`��J��Şk3��N�������;�.�,[�\7v�f]~����e��ʕk����[
HلR�M(qi8�O�R6;}�s9<�F~��w-��u��Jy��hY�����߼u[~�3�/�`�j=�1WD�]��ZH�����Ts�}E��U�-1�œv���P���<e���P��00OAJ��$��'�)��ҒK��/<1�O�ͩ�qG�L�:}�zcN��-`6�b4�Xz���hҐc9۟�'ۖ�w~S�WnKCo-��t���u�4��Fbt������G��O�k2�u~��~�"�k2�p�\��֬!�&Sx������u]����r�[:�z��Fڦ�%����6�f0fq��,�>̛� 3캛���R�D�q"#u"K�͕���|�$/�[������s��yf�ॽ��]*j���Ե�M�� �鮷	����逷z�DK��jه��d[_`��Y�x�A�9�����˅�DLS�z�9�����ݩ��u�� @������^�h��٩/��)��1ȴOF�6���^S�>��I�Ve;�Ǯ� k;��AZ�˹YN *a ��X0�gM�s&�j���-Jk'�e)�©
	f�Tj����c�k��J�<�;V��6�F�G$���ɧ�}(��we}�EY���W�b�ҟ�vdm����� Қue2���}$�������l������:^s����rrx"gg'�Wo�����/k�s�-ݢ��ufe�Ajk�\��\������vT(���s��ז{2��e1�9���â_�������@�#f�Id�PDc�Q6 ��1���>H�a:;;�ޑ��C���T6�v�g:�Τ	Ob��ɱ��#w��j!�є�~�tnME�<�q������cUAy���w�����6�%?z��8�C{84  ��IDAT��f������@<63�4j�-, �\���!���ǀ�����JY枆H`�p�3Vss�MS�R�Ӻ #V��!@����ޭ�� ��@�qMؽY�='^���{*��Yk+)c�`��u���3;�B���r�޻R6���{[��n��ݔ:4&;7��t3܋�2y����?����[_ߕ?���˱Q�Q���O�Фw^|Q�ֻ4�pf)R�Ì�=1{��u�R`��Z@H�A��2�~%�#��K �P��}��w�g�"�g�V��!�a��R�T=�V��{��R
vdĥ�JK'�ѣٸr.�g:�r�����ns�ƺ��d(ҍ�l�[[�<<�\�7�44�˽/ʯ ����0��q��_y�g�%�����rZ�.���{V�vV]�rYE�^����/�4�!����k�pOA͆��@{'���@Q.��R��$:!��-�k�<��)�Y#�0rpG��g#_Q/����
!*��]pgO*o��0��B;���5M�[�	@����0����_X%�4El��;T&�ϧ����j�E%�Wx�W=B S����������=Y�>���%G�!�[����M/K��ސ����?�B���$s��:]�����t4�^<��a��˷n���+���Y☬�T�C"6�ZҒZ� 	�8�/��Ac�ܣاsd%k����oR�ؔÙcH,�#�f%��>Z�D2�8/����\zE����p�甼�� �z��^6�%��eSz�/ꝷߒ���?�V��xQ��6�+��-��x��#��vrR��ѐ��@�D�0ٗ7�����TEpQ��W#��n��>#/5�d��������{k��}:(��f𱰊҉_��,wz�@%C��D���~˝�v@S��)��7� eZp��X�z?O�W�;��wPkb��!К�Yh9��d�NW.����mL>������A`��x*��Y�h���+�Y�L.���;RoL�6�m�7���b�)�u` BY�x.k�8�eOk�?�yU�}-al�������@:W��0
�z�O���L����%��LS�S	���y�)K�3�8�͒{��NO�&?4сC=�	6�(4��˭%���֣����ymW���!�Z��ST�ʐ/���\��������_�A����BN��������-Xf ��6`%���W
D���0�&@��Z�7�җ���Hô�Y�`L˨/���qu�u��YD�:sgey3^�E�㐼âI�r���7�Ig87bo[O	����
�A���XC���2���Ő�r��Y���x$g�}��s��@$�၁1�Qk�Y��%�
�y��l�2���v >Q�&�kXa��w4/:5]��W�p��>c 6���gBs��W%�:v�)����^�����˸�1�n ��c�"��A�J�r�_y�����}[�ԩ��=ZШ'�>��5�1 �8Z����T�)��9�u48EH�e)&����6@]����F��u�\y�H'I�#��w�Cpx2म7dW:99��޵Dh�rs�kzn�^@�"~�-r���䜘����]P���e\�z���$8Pm�ł
݋��(��4z������0.{��nR�Lc0� ���3�a�Ŝ��K��J�D=8;2��np.�A��K�f�� u�I��(�����g]������p�@�xHZG*����Nμ�� �eN�P>�ӵ�w45-�c��&5`����c.ع��0��`�¼?ưf�pva=�����������,��<� GGg������;���c�v��_x�r[��.��{�r~v&��M��0�f#	8��b/N�K��_p��8,W��C�}U�!�����]o��������rn �ȝ���9��"�c`4�H�ؑ�tB�®�*;SB��	!�-�3���!�j-KR��KFT�*���O��ݱ4��[��ʀ�Y"3}|Iφ~�X�Ҹ2HPFN�nWv�[&<]���<�1f$��N�nm�@��f��-�tN�&l�zxZLB3��j_����n�I�T,��_q��Q�%�"P��1Җ����w%$�H<�e��*C�p�X@3�Z
�Ԙǰ~���dޔ5\ѳ�=��^N�9�%�`54��Dx S��j�FDbcs=4=���u��ۖ�ӹ�
3��?����_���,R�s�?��֚�����]��^����X�Qs7h��~��u���:G�=�Oc�����������!`��L�t�ݘ~>vz�"~�U����g&Qa]@�Y�+�p�q	�sE��Gah?��l^�#Z3���v��؋�Љo��z� S�LB�p�O^��E^�cƞ�(�YOb_����%�y�gn�b&�`TS��ר0����{>`x�d�c���O��n�KEt�g��O��\�ƺ[�A_%��-a�ⰠC�VxE����b)�,��͝��Y"��s+|���gG�UY,���Q��VV�X��(���nN�#�Ʈ�ht4LP7,�䭷o�h��"���������JHD�7���4�(��2sss[_|,�|$)��P#ύ"~���Ҏzy�G+h�'���<���Ŧ �v���ʹ�e�9����������׺��;�.ιS�c���-�"����Tc隴�`�2BSp�l�&�IL�%6���E[\���bp��e�V�&e)��-�,=�v N�}3�ƙ�s�P��3u��wV��FyG�Op^DW��۸����� d�8���I���'��'`����l���w��Z1ȫL��h��NY=���&���>�6|����Q�>y.�O��U��J��j��p�P�aGJo|��Y�;�3�a��o�nV�����Ti�؄��Ra�00)�Ƥ��%�M�����r��������w;���7ų�uO� ����| |�N�YL�A�K�,=�2�
L8L����li�kD��&�. ���Wʌ˩x�(��g?�=��
�b��S��d��=<ph�dj��=��ʫwvm���ml��L}�ar`�`@�����Ԡ��&s
��[���&�C)�c)4�Fl���'ɍz��+�8�_�޵#��J��#3�EP�ĩ%�5ppW�CI/w�����,D ��9@WjT��]��.n;:W*=f��$g[vCB��t � ��l��b!�f��X����1�!�cm��4K*��(3	]�!�*]���3r��5���7���
�>��#�M\6��L,���q0L
�״<��/=�`�Ӷ^*�b��Z=:�_$��Y��tz�ך����'ku0��5 �k�[ǘ䦢T��>k��V[��Oޗ�j4n����jq�7|�#�! ��YL�.rI�s��*�@��ٶs��F���"�8eإ|0���\Y��(��hH�h,c�p��������F`�I��@$��m�Ι�F�%��\d�.�~_I�x+텧!I�Qh¡�TNh\��U`�����JSs)H�����ci�'�uc����IG��5jb4�3��%�і�ޖ�xbB,i�	�pQ����_I �	�D�{sU!���� a	�W��+%P����}K��Lo�4&n=P�
�)V��L�x}
obe#��<q)8�@�E.�#�9�k�Y�R��˰�G��'��L�&b��h�Ԟ��0�����b�9�jQ�����Ai�rO�2(v�H�&[��(�������ǵ��-��WqjIꘕ�z5��+��e��&��=�h`l�a.���s%!߶�M�[��L�A�;���2 Qt���8(�ۑ��;��{�-J�)��@>�Ahǲ���!ȹ������_��l�_�GG3�5��b^Y_��:L�%��X�x�*QM1�~/wy���X]Ș��������X�.Z��n�ai$�W�ܔ��lfo�j��Y�K͸���b^��)�=K1�x���5uncZ�d>�-��`�.lחm��r,�F�Ŭ@$���C(В\�f��ɂ0U�<~�//��m�/���N��S�?җ9�itl%�x�wtkn�^�=��6T�ʌ��k�h���MN1$����ǆ��].�=�de�L�5t<#�s[()�;bcѶWoތ}�����%bm���4�8�[Yө��
�<0-y肈"�<��$��T�yy0�A�%T)��*!a�����*W�
xPC��k�\�2D_�̋��>s��Mz�:ϗ"N���ê([�g�"�d�Y��v����~�R�<�˹{�I��_��.��>�X^�sS�?ߗ��u9��Go$OT�����}�s)u��V6��(�ƫrwd-V�E�p�h$�'�&̖p6t����ly��,-2� � ~6_D�=��Q�	j��{G�1?KBU���e��J�$�w�a2F֩�(�\ �Y�k�^������B]D�͋���u��4|s.���Ӗ-��bS,�i�4�&�b6��11���<�<�3�_��esG_\[zWK��Ϥ3�ʽ����r��.cuz:�����X9��`�B��(�R�ҕ��Eae6�e�`�0�����ز��9W��yiހ�wۜ�2[L(�
���O��Y�ª%���a���X���e��D�x�lc-х1��L*L"�'�W�S�8F̙$���Qp�}�G���y�5�.���z<A_^���ܬ�*�}.�rm���7r@įxr������G.RՌ�ڛ���\��U�@d��~����*l�䓏>  dGu�3$���w�6����qEV��Xfp6ָ�HNޗ�����h�ͷ~�X����Sn7��������Y���SW� 2=��Af޼[��a�猇"�'�ۓ:�~FbS�@�qg�t�R�h�sn���7im��j��/T��	%͎�7`�J�/Z���ԵK/uanE�B ���d�Ф������WS�.�� y~��zO  �]�͖\��ILL��_�z����W��hLO �`A݋�p���#�68��q�ò��	�Uļ�BIa����Fj��y�3I"O��'���S���H�%������"SbdZ�Z�W{|iY�#�4���9�6kb&3�$��@��������i�P(/�x�`t.V�S-5DC<_0��HQrK8J,���15a,��rU!#�'4�I���2���a�v�K�-�dx�]5֞��oT9�RV�!��bXy�@�d��1`>��e`RM�3�я~,�7ߐ��������Qn޼id�z��!wA���Ii�������[r� �+�ܸ����CB�����/H&R��k,���c�:�>��_ʴ�Ixe華�m��'��k4u��X�m/؁8�lN����L�KT.n��nM&�.��NN�&�\������s�&�t����ٻzk��[�a� ���ރ�@�zC���85���jZT�*Ɂ1Q��q}��z�-�'kzo��>�z`��O5�k���1�u�{r؏Q{8�}�GD�=����6;���bmj��!�h_���c��d�F�bw�,��B%��
�Œ���r���`׀#tP0�Ab�&d��,�"�ҥ'\�[P�`ވ2��,�c�Y�*�l����^�S�-�!��Zr��0���$[sĎh$&�3J�aK��b���j�,�[���pwӜ�����/1�s�jF���\J�K�K�]�uk��ܗn��Up�=���W���8TC�_�S��7�ȼ2�AK{�`μb�I~;��LT�¨���j�5}��e/W�}0�s���k��@O;�.'_ʭ�~M�?:����Pnl�Y�B#�9�:��Py>�Ȯ�Y���:ʢ�d>z$����Ϥ�qS^yiKF�C4^tSM0����C(��~�!K����c&�Ӟ�4F�G,2<��	��7ֶ�*c�4�����u��l��L���HC~��U���btx�� S5�.�3]�`�f2m�����/(���bJ�N�K��[���w��茽���Wz�����n�S��M:����:Q�"vg�Q��dtIiQ��xd%.��z�PϚ5�\dM���C5��H^x�©�R!k�m5D�	9�&I����� ��ƭ0A�� ��V�!�M���C5vQ*gŦ��,><ˋ��x�U�:4د����)�d#����6y�<$�tn�xl%�;iMV4��f]G�t�U%Q[K�\���%U��3�B:n��)�턦��J�b^C�`0b? ��o���tMC2pU��}�C�,�����������Ć�t� ���Z�;6>ؔ�-W��4�Dvt~%��01!��KdeN���e�!��~�w~Kn�rW>��syt���ژ@�f�"�<���.�N&}������>�B=�V-����Pz/Oۯ�l�',7������(�RW��BK��[�q�����kNd�;��|(���N���N��xI�}��:Չ�O�>���>�{��kꅴ����%�N5�0���ŋ��>��t�	8=�;t7X�8�a80Эr%��w�t<"]���D��LE,��\1��L�j ֶ%����tzk�� $�qHg��Ѡ�f#i�aB_K���
���_�9�nc�{A)3N�2�����8���{�������zG��3y�$c�)Ш �ip���S�.k�}�(���MT�3c9FaHY�6L]����uHZ7��l�Ͻ0j�� �A
}*j[.GX9Y�3�M,�����/g�T�eG-�^@�=���C�W�?��[��!'���R�u��
+��\N�Є���֘�-�GX�����=�X�^XY�,Amy���%
#�x�e�,��1��1D''4V�W�h[��E�m�r��K���E^�Y���Ihp��I�h\�/���iw,atvr*�Ǻн�,R����a��0MYi<�e���n��g� ���6=����N�V���!�<Н���3��ڏ~./޹�8.nO���$�Ȋ�e�`�Ȥ��ԅ>�b6��3�瞀��m����]�� �Ŝz�ꮀ?`�j��F�\b�1�������(��ce����x�'��)*=`E&eX�]�HL�EGh��v�*�$V�Qӓ�	6/�)���2�W���`l�W�A���0�C���sZ3���Z3ٺrE=����sK��)���B��Q�ca�A�ű;![؄�Z�����ʺ˶����
��/ZxE�b���jZ%[Df6A��c6������ܭf?Hb	�Ռ����R��p��Q�Hƙ:4��IU7��8�Gļ�j�p���a��Nź-�������B	
O|f�<��ᆁIKo�.W�
����r�\��eE3���i�h�m�s���*I���p��(���#��qQ݂�>���k��{�������&��e�u�>�����Ǐ6�232����b�*�beK2e�6�4������S�-�xd[H�DY$M�DBE��������>2����o^s�=>k����Y�+3��޻��sv���kJ=Z�����V�q���m{���������ݺɖv��9����n�[�W5����v�����v��X0���O�y��rQ7pK��p�:)��ɳzPj�|~qj��LE�~�9�5?������uv�ڑݼ�o��Oj���F�v�zԚ7Oz�M��b��5[�w^�'����xY߰gC3�UݘO����֑M�mV�՛o��!���?!���ݩ��&[h�>�^���� _և���>o�+Au�[7LM�06~��
�G��}�n=���s����j
Q��֞=������M����s�ھk[�@-O��N%�<8��;?{�qq'�}��Ckjd��7�nG/��}��~�����"�j�v���^��ˬiO�-F�]��xඡ~A�"���o\TG��t�����ù�͏��J��ا�4ԥ-^�����#���>dIri�=t+�wQ<�X}JTܰ�9 /#�"���|��@��bd�4͎�(S�E�Y�b����1`X�e��i&�핇 ����jZ�dpeC��J�@iq��c��&��&�a���ƙ�q�[W��6ʣ���SEP}�ƭz�)�/�E�PuM���T�ok�H��u��.�H8-|�C��P8�󺏐R��Y�Q�̫�^������G��r��V���uOkd���َ^��������c����:���+ ��[SC�[���;:�a7�nш�/�WϹ��v�E�v��w�|�n��En���k� 8���}{v�Ȏjʲw��铏�!޳{/�S���=~P�~=�/[�w�Y50�G��s�#��\^�lk���0�a��H��v�%�ۖ6Ƴ��?�g	���c�_�C\��e�K��=���5Ӧo1:؞�&��0���j�Հt�s�^˳��fvvf��ݴ�o�Ծx���=��۞ZY?�����%[�hǏ?�[_y��������[vp�����ٽ7�`����Ӛ����_���{�6*�f'���l�FC�6�]�������J2��-{�ŗ�z@��&��>ˑ��H�]@�j��'�9҃��D��U��)���r68/{U��Ro�P��IZ>�&c�} f\iym��`����!��a�T�?y�k�>��9���T5��� �G�1DQ�F�%�7�D4v�f��[R���%���(�OhL�� "V�FViHw�d(���g{o6���ڲ�� �h��ԫtM\lq�xZջ��N3�Y� RnC@4&���v�k(@���[שt{�s�:�g�s?������߶�?���jhN�-�U�W���O���ް���Ո�n�zpv>�E�<�)��5��y=@��<����%p\��F�vؽk�/����ڗO�Z[�gv���vPګ�B5T��9�k�_��F*ˇ�ح�{��Գ��n:��sݮ��_s�쨽n���>���|�W�j��rh5{��ގ-��Hi�.�*���li����m=�F���"����b݃�=�k��mv���_��wl�-�<��'g�rW�19�����O�!�ߩi�'Ղϫ;���:$�������zm'�\<����#螢���P�3��jnZ���ӻf;ԥ|���uG=�fulg���{hOm���e�n��5��s�"؈�]*ԅ�m���"Gr��+���kڤѵ(��^��)*�1���YY��5o!M�ZI�{��:�TmhSt}CŃ�a�x��4P��H������G���T�4������� ���!��oA�*�Y�8�M"s���)i��m�%X����b:���5��v` �Z�W6xT��C;� 0ٝ�9Re%���c�E�5#��z:�k�1b�;M:�P�0Fަ*S��]4ݻ�2��2Z����w샏?����R�~.9��K�5o����7?��z��vn���ß�؞>~�����?���G�����~Z�{5�_��y����>����(����Z��=��
���ل����߫�򬆙;�}t^�Ϛ�<~����6}rA���?�����S�`���ʖJ������������Y��h.{Rÿ��#;;9��~c�=��j�?}bG7n�����nk�O߮�{n�}���ql��3n�/�(��ީ�1!s����>��F9;;v����?�������� =�����)�r���E�Ok�o�?��]��o��{�O/)����9K�ON���9���xj�'�H�y_juhgOQ�ص�O>����=�Y�t��xNgu�&��Ow��˯_V2��f��#�װx�����x����Fg��*�\;�y1x��IՇ(���V#��t���(@4Мٱ�X� �p!�϶pd�����G�k0hfK�ޟ (u2z�M�y/�?ל@�WG��#"U���O�.��^Ո��<����W���9�I�2Lr����R>�g�Y�a5R�%�1&��z�)��©h�`;2������A��0�-}B�7������8D/�t����wo� �?{��5�5g�#հ����K_����{��U/�={��95?I�<=��Y�E5��O�������zɳ�쑇�yr��v������H�|��E�6�N/�l��E�@�������Ӛr��͜������v�����_ӟ�<�QpV�~��Y�n
����������gu�q $ϻ�m�~�g�9Z\���o�5�>��o�?$�m��tn�|�->��=��������5'�����7m��vv��F#H�ۛݬ��>�z��9��=�����uM��uMw&ŶS�N�z�wj$���ϟ�^��~�����i��5Ҙ��bVc�>�g5�ګi��޶=����K]�[Gՠ,��?�������|�Z����C�uR�K���@ �jr��b��JƂ������$�J.@i��%?�ز��A��.P�m��@g������f�{gJ��������c�!�dE�Ib�9(�3-�A6V��)�w�c�����Wf�L^[����ϱ�b:<�iT��0��TD�d�,iL������3���K�r�����|�6�Y�
ed��GyM�t=���g� �Q�fp6��+~���8�#ܭ���{�����g?�}d[�e�|��8dۺu��~�o�z�e���v��l���v0Kv��)�|�f�3&(V/���G)^��������=;�������XKTK�@a�1��BeH ��<������4��Q�\��~�4�?���A5X�vf��$N_�2����q���$?�_)�ݚdF(��z�[;?9�weU��)��h�2�A5�+� �2��5[vX�H�?��o��+���˽r�UN�z��?���uM_ ܲ��C�_��yݼ��ޢ
T�(���GQ`h-�Y-ˤ�뚲M��`~h��U�xRS��}��ͷ�!�n�?���}�%�D�%�ը��]�(Q����U�+̻�LɎ�xx]E���C�Bg/��L�N�.���kc�(�oy_�	Q��WD3��0�g���C<��״������j��F~���u/f�8-�H�{x��
� �!�J�H�D%y��>1�"��(�0����IQI�����j���+�O�?��+	ܤ��i���W�>s|GeM�=�:�d>�2Y� �����d~d?���?�GOO��}����6��J�ۏ�я�kݓ�lu���LQn�j�w�J��G��Q���/�tU����n����]۱�����A�`s۹v�z�zP?�����^���58��] ��/��]r2�%��@x<��W�}��2�[��rA������u�_���nݼU��Ք���ݻ����V5����ӧ����9]S�3j��ޝ[/���4��Q��xVӌ�/|�^�S�L[�Y�.;������;������vX><�S��y��s�]���m�7w�O���70�f�ބ����ᑭ'[��f��1���<��˲����ЯY��&w^���n=���}�A5�3{X7�i5��݆:�}5��.��������߰kո|�˟���k�7]���H��b��{�9�:�j�q�MR�qhȳh���
:�+S�lu	J���������0m6<۵�]d1�����D �p���V�1�T	@���	�����k�?�p37!ۗ�d�4��������H�R��;e$J������&�i��?1S�՜�w�q\���4N�nI���c�s$׶3,��J ����.S��bZWT���9��64�Xc�\8T�Ab枠�@i�'�O��;/�k��Z��S��j��ٙ����_���Ţ>���/ذ_�/}��/ڲ�ٝ�۝o�q��gu��V/z����۽/���l��-.���E��{/�l�o�k�p���E�=9��^~�~�wۖ5,��׬�����o?���������3n��[�s�����ն�g�����ݷ�g��������k�`��?��޷�|����|`_{�Wl��]{��g�������v��g�>����q'�/���������=x�=��>�׿�s�����i�^y��?}ˮ]�I����-;��d��?�7�����߲Ã{��G�n�G��?�#��7���o��oڏ>�c��~�>�da������7���oo���޾��_��ra��ݳ��C��������~l�������E;;�����S����[��k'�b���_��~`o��]�|lg��֝�v���n�}Ŷv���w޷��'�״��ڞ��կ���j��<�k{��8�@�svi�H��=_w���=t��lH܅��Y�#��۵5��@������6<�*v�(:.��ئ��f�`��A��X��Jh�O���6�_@9
�?J��En��3�ٙ�}/ؖ5���-�^	ܗ�TQ�! �t�TQ���5x$P�����F㩆�xy������DO�ux�J/�;�f�>�m�j#Д�MSֲ3QE�*�h=��h�0���?���S���F�2�O�c�?sptd��x�_������{�ߞ~��m�ʰ�i�,��U4I�2�nn��Սpkˮ���t� �^}`o��Y~z�܄�?��5ǿ_�<���]R���ko�[���]��_�E�>��@�ž�K������c����ر]3��o�<�����{54���iڵ��w������k4�������o��m+[��'?��?b�á-�k��Gj/����o�����i?}�c�>��7��޶A�>]��^��ɟ���o��ޛ�����/O촆�'�g����ؾ����<_��j�n~ƞ��`��}߆W�qX���ĞU#���G��[ߧ�ٓ�\�}�G��{QS	�N�уs�n�o�5������}�����??f.��w߲?��>^�<����[?���	 �����5�8gCխ�wY.����69�� �TC����m��	����EWb?x�R�����N��r����co
K��Ė~�_и^�>ɩn`�j"2R(1��@8��L\�e�S�D^����;���D�H�tu�ڱ��r�:tk4�X��a��y8o=+4�����\����C�z7<{Kŭ5:���`�,�3k�J�J�3t:�����vl�#m��#I�������X�G��l�И��Ө-(���Z�����Mj豺P9�B:Q~Ӳ��Qj�&�bv��`� Hܞ��������W_���L�b]�W��J�_�����G߶��wj�q�ֳ8�E!��P�iC?��N�r��;�~�����7���������_~�_���c~紆�� ������`i�m��a:?`��®����?�}[l���x�1V��o�/4Vm��>z����ϞU�qhO�C�{������M[������\���s����A(���>�l���W�y�v=P/��xr���5u�u���<�U����O짟<��|�K�O~���iˉ�������v^7$<�{��������k����ũ�����?{f�o^��|�����o��rq�P���?���B�@�><BE�]�v�v���=��{�Wlo�
<�����-����v��}������]�~t��}��k��Ė�FX�09�A��
+�u������A!��!9����#�Ͽ�D[����:� �r���L��6�����ȫ
Q��	�.z��?>����Ϟ�6�')[�I�ް��-�[�3t8)�CæI���� `?j�a�M3c2���#_�`#�R�:˪�#B�G!�C��^�MS���(Q�v�¸��jDKBVO+`)�;�2"��F�+Z�ָ�\E?�F@b1K�#�^Y�x@I2As��9+l�B��*����}��7l]7ⳡ�۶�5v�����or�֤�b��n� �=��=�9i��;�`\?�av���f��g��_��->z�vla�5ʘ�=��^;����������~f�}�̿t��g��żV��/q���G�j�����.V���_�a_��|�j�� `�vfs[��f�	�<�g?>>�����9 �^�}���P�	��^�n�/�/�}�>�)�!�_��-//h巼T�6k�y��g�5¸q�==9�{/�d���A=P���B*F�,S�{w���F��\�A�U��u�Ofv�\�+�*S��;��e�찦d����u�a'g)1�W#@�-r�䢎�F鈕4�z�G�B�+�$oV�J�x0ս����iX���=pLH#��da�tX�+%:�V����D�%9B�`��0$�ʠ,�ƹF*���8�T�.��%|,]�LQ��T��y��ѹ)n���F�"r�">���"26��B��Ml3^�؈���
�m،���h��1���LJY�u\�ϱQ�QJ�ֆ+��iK�H"
%�G`���j���e[��oh�qD{1r��]�,�_��������k��޵�م�M{�qt�N��)�g���;�	S���Q5+�~oԐvR��ç*gA���ݯ�Ξ`��U�vKy�F3�����^\��C�5�7��!�O�k��[���d%��]���]olf?��;�v�y)*&�w�1/��۱'>�^��V���h��'��j�����X|��-z��'O��uN���=V(����zMոlo�����9H5��O���q@������d*�,^�8�D�u�Fvٝ�,�a��.�i]��������<���ޘ�h���.����s\$�^�d>qť��hs�G��xĿ7iDً�1��B���˕ʑus��\�qC�;�$�/�.����;@�w��l���"�-�loh<�$ul��8'w��07;0�u]����!?lD���& C�^ښ���FU�Ƀ�x��)!��z��gٷx�$/S�	��A�1�U�[����9���SxĔe3���`�ᰦ`��P�2'c%��G�29#s3���(ELØ��p�q�z�9� ���ҚԷ{��m˻Kl;ƨ������[^ֿ��zf<�U:�g�6Kk=B�z�� }��c�n����F��ݪY�ؐgv��ω������=!�S�څ
SWn�w����ݙB��輟�o*���Ŗ(3C>�Zͭz(�(�����~X�z�E9�k2?�ơ�}��2�u_�j��t6�Ϣ�������nZ���A�j�^t�S��j�����u{�RxsPs%>����	�!p�h�Z�(
�p�$
��ن� �尚w�W/�����fy�qMK���|��>GI�j��Ԣ�<����7�� ��&:m��-��#6j�?v�<�	��h��8�ܨ!e�??��Lqo/�|����:*:�:�9��k����vV[R��$�ّ�TKz��_�R8{�%�@�F)N��OQ^��j���Qh@�Z�Ē���}�:��q-�,�M]cV�tj�6�� �3N���4��u�����|��+>���?��g�%)�+G�6C��T���]���IL�,��S�p�݃7�vqv�z�5�F.Z=����+��W2&2U��/\��e+v���Þ�M<%E4�Pe:�!᪙@Pu�uh�<֚����J(/.jx���e���]�?�lZ��i}���KOj�|h���3z!��Rc��Z;��5����jT�\84�H3����V����wC5�CN���D�aj�t�.��`66J������d&����>9GE���v��h����7Ѽ�f���a����f�������-N@�Ԅ`<�,;-�8����@���qW���2o96
a�Ʊ%bEz����*�8*Ό�sD#�Vmmv�b���	?|�M�^��/�VD7h�IJ�����U�$�^�=y�u��q���Oc�2*=����(���Ք���S��A��
b��� @�����=��=�#=0�6�q(�?� 톷04nJ�Ϳ��LF��G��D��?o�E�]�67Q^̤֩y�ð�q���ƥUi����n=��X����
�u���2t�s�5olT�<���5u'�����z��C���>�	5��^�dlY@�����!�K�*q�:�ug�T�pg�r֮���F�ߚ�L1�����p�9��zj�/������K���A��u�,���+V[�L� U?���c�nv�Ĉ�킫0\���H�ڙ7�ۏ�O�`�P�:T�f���<�Q#P;�G�w���y@�P���/�-��d�B�3iw��.�g�`[�m�U0TTP.�7�j��t�����bN�*e!/�"@榭F|uN�o��������؃���%��#����G]�>I��3���_E����3ښWJu��r�|�>�e)�}iR�O�6��E����[ı(��ل���b�Q|ȱI��0ph��$��n{�fW�'�۩�嚯(?����\b��ަΠi��p�;[tTo�9N����� zj\�fZ�Y�i����o�9LZæ8y�b4>a�i�{��ڕ��OR������uw3'���wj�?�h@BBc�ꛦ>�H}ﭶ��\b-4�u�-�,o���0N�9�N��ķ5?P~Ǻ���Ԙ.H�-l}�L���9�n�U��e��ŀ@/��#</�pf
��g��҈�UO�>�n��N7q`�%�U�u��c�1#���z�jtE5{��{��\��ꉞ?f��sV"��)�0���c�}�=;>�t!2�<���ț�C�Wu��4hb���Y(� $|��~}�',�!���+/�����a�X��6ӣ���O�x� ��ΦdE�j� б�Y����R�R�և����.�j�!�g�?������B|�#���O��HCC�F��0�
0Oe���J�{�/*bp5eXN��q��*j_�(��04�{sz)��
�IV>90����')���K3>���>Htq�A�`�aM3H��J����>���J�x�	:4.Þ]~_���4b=��)v�Djr�覵�u"�\i�������m�;P�g^���$�H��-T��|v�)L�Ȯ&oI�
y����y�<�CA(��j�[���"u���w�X,�sS����2R�>ĵ��L���ad���"#TZ�T�]/V�O8ܵz֋%�hv�f�����&Ld	1�j�K�w���^�aDi�(<"�Y!;J_r�uqvL�j �6��r��oխ�����5;�U�fت����9M	^��&����J3Z��,@ж�mfI�1��[\.5f�����e�L���Uk<k�G��ǉF�����h�Gg���%²	�pr�/���>DjS�n(V1tWތ5iӖ���l�N�a����Dh�CP���7�c�5���;[�Pd�b��e��QE%9����vK�!I&�hc��ꂟ���/h�T�J?�T�����<�6rEK����3�nE~���jtZ#A�;��6�7L��z�}zvy�q-:`�>6@���1���
�	�4>x�#������աA��>@�Q��݆P1M�ֽ�Oj ��#a��""�;gU�x�Z6V8F�,<o4-���k�k_-�s ��Fn,�G����S�#X���Z���dUBb74�ׁ�'K"���,�0(����~�*7I�~�"O��&Ʒ �Y�f��B�����1ql��C,�$�i^O��U�(�‖��������l#�Nmo�͗aq/���Z'������#�j�>� �{w����*j��{�g@R�'Q�B�.RkD�������	��t<:��tez���W5�;�gR�6:�x!�@�0�U���;#S{T��j�*ĳ42��j���@�r�ة�'���u|��G]S�N�,�s
�dP�mAU�u�@AO�����.5��,�h�WĤ��-�ӱ�vpD�qH(��j89M�r{��m������dDǕ!���b��
��N7~oJ�?��T�����Q;qE����̊��D䡇�RՇ��R�B���f��-EK�kb��JA0|�A��}�R��۱鱮���k�
�{H^6*A-.2���}x� D�G����8.})^�����^�=T�Ɇ����&�+�'��S�q�H�5��u1ѫs���T������@��ǖ��Kʏ�$'�� ��{�K�8ML�7�5<l��f���Nk�C�œ�B���i�M� b�"$��O+�saJ��{J�Dx�� ��d�N5ю7�#-#s�p�)u+(c���,B��@N�ĲP�8�J^q�2*kq�G��E�񦫁s,�Kӊ��� ��Kcij��AVF͋�z<��N]Xl:�ߋ��v�DAMƶas�|<T�a>�8Qd-o���]��'P_%���xm��dixp/�0`D%�FJD��8(��f��6�]���#�W ��oq���$� ��8g����N>:N������ɀ�St�@�x�l:c\%�����E����wj�Vi��p7����k�KBGeq�}�1���N�`��̹!��5D�����x�e�
�}��Z\�h\�X�U2�3�s�{C��l�e�Bg�4`<����%�S %]V���	�ك�"x_�V�֢X��M���¾�q_D�Ӑ��Q ��N٩��Tq��(��9";^0�+e^4Wk���i��m�Ŗ�I079a�hY����h���O�˭��L&����Ŭ���Q7��)\S(�YC�Fzo�Nn���B�Di ��<H ��;߄���l�|o��dx��M3	�1\Q��4𠠌(����ʱgIy�
�����D��N����XE*�����k靺�R�{�(��h/J��7��+�]����
�'��{X���t���?p�ɋ7r�a8&5�M�wMm������r��8�-E�OVm��Њ'���.]���l�2�;�p�vC��c���F���7�(���>wO�@�Y�̻�a��Z6�n=�
�����kV��j(pV�ʰ�s;���}(�A�\���,�9;��Y [AI���(�o� (
�e4X�.0PQ�27X��O>��脢���FV:���#.���it0p�����^-�ko�d*�xfY#��`���,Vd|�Z�KjMf�Q B�� Ք䉵�=2��]ź�@��ƫEQ�-�B�|[�(1O9�YO��}A�w#���=�o���Q���Wx���a��� ��_��"fD�ϊQs:�q'"Sm���C������7���\/�X�Y ܦN���-B|��0��Fsl�z��SL��8x�@p�c��Q�1��],/F¢���!�I�
6���)��B���+��A��{��z���E���>�3���C �D�5g!EE�:_�a�8�Ѭ���3��s�
D����R {�f<R�6Hޏ`bc��)�.kMd�� m��6krT��l�jJ���"�-��/Z�;�?Y��F�r�����Z?����}����R����^F�Y��U!�FbR�VLP��Wxg'�����[�}N�B�AD��VL�O9�gѧ�QE�S^���I��tPX��1$���+�+u=
�j\ٯh��J��F9����5)�����>��k#��1�`��$6V��H(�D:�I(�G����>Omp��:8aC�K ���R��5����Ѱ_x��²G����^�Gf�~x���X¬�4��x�p:�P�r\�YĔ�(�� ��WE<�䓒D\��$�. �k�����}`iS����!��fI�R�E>���O?#�Tɑh'b�׺����Gc���ڳ��k�6i.���.,�W|�D/���(A%��fQ�C�:3M�dd2xD�6>��&/�jt�COPu=FN漃���S\Fak|��r�Ӟj���Fry�_����{@^n�on���½�$�R�
{�F�#�boP�ׯ3q�H��\��6T�:/��V��<���"ꀦ�O�7X���C�u�Z���!�WB��R �~ ��|��y������4��X���L(�1Eȏ��AB-i���6�����7-'W�q�x�K�e��ǁ�������K��z��s�}�5O��}�
���n� �h��c�Gϥߔ�ǘǇ�d1�-�F��K���kW$�����Z��2R�k�LTjt7k��)x(�bn4J�aH�ԍR�u�*q03I�qZ���+S�ږQu?��2����+�H�L<l��I��K���]�����ӳ�4�t,��:Qy�d�Ʊ����S3Ifd��3�����=U<8� ����W�qF`��=�f(=i�<K�O��"�4U;�C|nh�.륞	�8�̓;��
���4�<�32�'	����9��!����.֯F����{N��v����p��q
�Pc �D�^�49�ҸRlEٙS{��f����-���~��p�HW�?�th�n�ao��;�(W=_!0�����wFk�B���A��+V�����dHe2X،��X(�0��5�i���$��@`�ΡlU�w�y6'7�4���,��lT�ñ�<x�d��!�P�2n�1?�(/�ݯ�(�7�9��H3^k}���x?�F�X4Ұ��BV�z\�	6T;U�1�w��6 ���x���]�������Kc��9(L9�^�[ t��xPI�?�O��k��vP�SX�!���P�̓1�}�h�4t�{��rSâ緳��Ĭ�< �Ŭ�?H�!� ]�	p4Y"ס�!��B�.֔�kw X�; ����Å�k��2�$1P
�(��C��q)S�Y�B:��=����:�H#"�.iW�"1�sa��Z� %��f0]K�9�]�'a��3��>���XSP�0}9��~�����jn�b��m!��Đ�}1�|�d>7�s���H@�^#�PC��K�Li�
�^M�c4��'v�9UDZиA��+�(����4^_��77�Z��y���J�@��r]�B��H�����e��Dt�8a���O�r�F�I�,�X�䩃��hI��f;:� i[CX�" ���W�s!� S�R�y�W��Ѱ�s��5��գ�L϶�����������K��N���� �\���'�B��#��	�U�����F2��Vg!��V�;eg��Ȟs��K���"�U|��ӄÛ��`^9q�dJC8��H1l&q�3�t1�+��,Jќ��恆��E���KڨhY(p���{���l#uD�˜�u����湘����w0q�yr��j�F����\)����&CR�,�L8���%9,D�-.V8�r�
0Y�*O`��{�O����C��9�w�4����l�)I�?�TY���`WҎ���{��6@墧� �Q��l���@�7ic��7� �́��w����֍H��1+	���)���
�A���Q�"����x���u���5���q=�: #m'{	d"������8Ѱ�m/³1��!���<� ѣ����U�����it�Zv�J�D�J��5@_��^?�:��
��幀fP� �SS�~�)W�4���Ĵ����Z�.Ԇ�2&N%�Cy�$��bN��T��[����N�h�x)�	)SYA(��������'ˋ���k��}��DN4����#�t);e�ݴ�K#��狨��ɐ&cO��Lㆺ��x��H�1Dt�Z����w�, �
;9�8D�^=L�%�� �` �����]�G���h�I#�>saA�P&~��N��Q!�\� ��@+�&|͊,�#���Le-�I ǆ�3
����*S���7�+�w�i;Fs�:������o�yH������]���RR�f�" ���#�F*]|tp�7:)=�ml�UerUhg�^-��#�Ȟ^dQ{�<ԡ�j��$�c��;sM1�sQ��n�~*�_�W�į~$)MV@��ȩ�(nm�@��7^r���bov�Ԣ���'��h5��'xd�T!���_��ҺZ�E��hd�2t�ٕ��Ok�����h�!D땀"�FV�a���4ޏkl6c9:���;�Gla:��5�aT�\�|[�뎓EǬ��T��{���6��Uh
��O���$�6��C���V�ZI��^7��Q�i���C� 4��^���ad�I-�D��V��ac�%4�"$�d���^ɨ�f���M���0VY�9�<��*|a͛q�����:m�(p&q���Fy���{c��H��1����f���T�"<*��!&���JP�`p�a/��f�mv�؅^6<_|�]u#ߐ��Fєм-ň9���p�<���5�����h�B���g�V��>@1 ���G�&l Li�6�A��d���.��يw��H�kx��Y՛ҏ aH��g;9�f|^��X."��2>x$�S��ZgEژs��s|��|ɫE0Z�p<���&N���_�F�����6�dQ0UU�fA;`���R��4��Cu1fb%Qve�c][�{�+��_����z}��R%ڷp�r���+ώ&�\�ӏL67"��mF�M �R�����&ϱ�w0���o) B	���1iHɨ4��Ϙ��lXٴ�"�HW��z�p<���Q�jmLbc�P�)��H�Jo�O-+���BL��1�u<C;���ʕٓ�:;b�^QDJ0�8�Q@��,�`���߃�0�A��I).,ث��s��c��$Iy�{{���{B����J�|/J����F�<q0��]�+�1�a��X��^����Ė����֊�0>���;�0Ҥ)��ɰ	��٫c�9�ȩי�pcj.�j\�����$RT �t��q�Ʊ�t?R�}E��z.b�?�ɸW��qH\�iZw�q	����q�U�}�]���HL�U��M�<`bH�)�(���������V���7��&�{�;e�t>����8ɞf$�X���?�QIp����Dy~z����"pMC�����}J6|c�UN-.�޸X�p76�t)�c3��.1��
H�W{���Ԏ!���d�;P� }`�=K�δ���V*��i�i�F�%־מ'�2@f�/j�5#��'��]Lj ��"/��^Q�H� p�	b�|@S��vׇ�&Jp
�t���h���_Ē"}t�8�+f6�i�:��yga�)�Wd(\�8�3H=�?S��{�9�2ޱJ��F]�da��W0��l����Ƞ�X�S��;I�8y&�fc�/�\��{Ϳ�hC7��%]��`yg)#ʰy�F�lri/�H�b����J��I�)�˴ӳ�޿O����h�\���u��"^�t6�V5;�e�)g������տ|�I��1vǍTOu�$���=�|m bG���PuX-֚�p�S�^u<�^|ő�6��*�wل���l�A��܌Tn�SF�OEi�xj�y,�n����� z�F9&#+���ܒ=j��`D����/j��P`�"˰ ���P����/b��I��f�Zz�!0��gb�Z���37��2��Ї��}>��DD�5;�[_8@-�!1��<+J�/�� 7Iv5Fl�n���z���ӎ�ʽq�ɔ�Ȃ��F�gE�eL)���A4�}9�����#ᱻ�S]n�Fq** 9�[kQI�|��v'��
�f���Q"��5l~�A6~�#
fh"�E�,{*�k��r�Z�i�=���u}%���[�v�̳���v�����nU#���X����RV�0��Z{������娱��ܢ��5���F𒨻�>���^����G�zw�k �h�M��
�y�fE�@�V�`��UpԨ��0��ƙd��0�ネ�KMö��G���&�e9hH,�K`lH1q�d�=�)����8�]}���o:����`B���8պn�&�'��x�߿{b��_��eq~�f�`��<�� �����>qa�"�i���=R�n�Zqe8�1�Ð�٤� O�A�xCK1d臢Yk�I��aJ��O�v줎[����"�^4EE�
�;u�z�(v�G�؜6��Њ Ѽ��H�+bR�J�\�3�"$�ϙ�! k���vP6D�4��+�e������{N^-D�T�,���͛�9�a��yHr��*b7;���)�'�m��I����b�?<=~j�{�,ڭG�1,�u�
�l�}OW詮�G�Bm�$c4�g��@�_\_Ș����6o�Fs}���e]!�D/�$odahi�eOJ(!#��G/����+0�C	
�|�D���ד��k( �Tc�FQ�u�ƨ�o�V�u�A)��n%ӽ�C]��^F��=����5�q>��LL��[�و^��I�ρ]����� �p����Y���q��HG#�\߃4z�T�3��fuw^��2��?�n�,zsq�3����y 7�(|s��h��	�A"Z�~%���|N�)`��Y�������I�Zp�^M�� ���H�2O�^�J���=��3$�5��I��阾O��f$S4&*��5P�\پ�i�k�����X�t'�?w�I���ť]ۿn�y۞/q�b���ZR��|Eo���&��YBiQrɬ��3��
f��npݫF`	Y'9�(&�W�,��9�yǉ����A��/O�-��p-Od<�AL�
���I)<3a���I��IQ�Bv���|�w��g6G��(�uf'���X''�]?��S09�i����FMsS��x�θ�Y�
ӯ1��`ݱxUxP+��P#Z�A*�F����Ez#��hzRŋ��"���H�I��N����0�	Ә�����Գ�vs��ш� ��i�<�{�m�7�Q��)U�9�|o�a W��Tkiq���%�P�� ��zȑЙ�,�A`�x�i+H�q�H�e�CHe`��u6x�7Ҿg�`9F��Ͼ$q�+����6�Y���Q�{PŇ)�̶�|^'{p�ݸv{e��r�PCcL��!�
�2d�C$s#�nQ�k�؛������� �n���"8��7��_ܴ��L]�f��ܥ��fᔲ{=�QEhOt^On�yH�gymD(��p J�X�S��I�U����T�������kVdC���7�V�� ��}q�7��)�V�Ӌb���=���K������Q���eE&�bSv}B��$Pp`���(Kv<S��s`M����td�ݦ*�8h��Q��QM� �)~p����j3!+:Z�L��4�%�û�:?�(�j�l�a�`� nʜ;��y%tGe ��e)\`2k���?=wlb�ރ�Ӗ+%�0� N��Jٳ��w�k��5o<���76~�9f��p��L����r��Ā�5�d����;���j��}�Wt����W]پ�K�`��=�8H��8�[5�|�.xW^\�,�9�9���#�b
Rv�� �p\(�N�2�� j"HyU�F���;����'�R�i�7��{SZn��4{��G"��ȓ� Μ�!F����ez�M�����sn����f��Z_,l�;%0F'���D||�z�͉�#����s.'�m�30C��K�B��c��Ё0�T�h���BX�Ѝ�~5��jD�2�����Dn�:�̈́�&�,A�����O%�v�-.�9����;ԭ�����I�^�;�3$�|�ڍH��InF���[9qM�]��&����s��`�Yc;��2����6T)c�>+W+>Oh$�h6�ȹ�CCS��?+���6
���y�.�6C|�;&P�Z�Zt��L���eg�hǽ�]�� EeO�� �ޱ��eS��]�\�[�8�|@���|�E��>��;�6�ݡ�e�$��S��nL�m�\X�aQ�m>��'j��%{�d����t�fJʭD*��)�=��P^���q���bF j�NX�̎��!3��ǃ�����l���E�<8GV9:F�fݦ>�`�8�!Dd|��l0��M�&k��E��� L��K��z���� �I�d�������K #K���,ґ�Ts� ?&���<��ә�ƃ�S��`T�zO������w���F
5�(�J�c����ǃ|��ӕ�|L�
f��=cd�L��y���È��4��-o"���^Dy2 r)V���dΕ�S�~	*(T,��+N����8!�D�d,��q#w'�I�'��~gR�[ȵV:���2�����>� ���g|�"�N� �����;x���&0	��tS1�T�"�!���|%D��h�N���������[p�rV>�	f4I������th'{dYE���eS;3�L7փ��A�	��oqk�{�br�Qs��m��$1Ս�"=hU5 zL�K�dO;���Eށ�W��B9�����F�0e��.`J��֛��>DvQ[8�y����˼	t�-�jZ�uϱq��x�U>LQ�;�&����RI���׹�Âe:x_�rf\`P��G4):`H݋R��/���-hH�5�IF*��s��N���:X��@�.��P>�lٲwٸ�kQ��h5��+���E�pv�����]._׸��@�Dǲ�w���؜�2 �H�F�p�.>�h����<7�/Z_h�Q�`��
6���RN���!�٠"8��ts%,i>��°�Pa��^��{#�e6߶��7l���T�,����fԔ��F����:�%(i�i@ bH����V-�,І7��F�\㔟�S�������8�y)/��!x�Y �0q��M+�4J�+�V�*Z��X zWI�ہ���b�NZ�1 �; wM�oH��/�1V(Y<RP�%"��B�M>�Ff�с+��s5e$��;�����
��(%�嘼aI��lH��ԯ�Ԗ�atl��#��t�o���Px�.�q1́�P�$�����x�����9ayi+��[����K~D>{iX�?c�g���d�ʦ�S�J����G���"}��=<T2O
� �l�<*�,�Ia�D(�ZuE���1���=��M`0�6��AE<��^�g����D#rl�o'.Z3p֭����F�1�$��1��g���
��^��B>AN�⭖�[׍�� [�������H��k����K*K|ʪm� &�8�O�*�jM�+	���Ɯ*J�l�"������0�wV-��b�2	e������������3Z������g?����{�E�����MY4�����P�rh�D9�&Ͻl%�
��97��XՖ��� �1{Q��rp��:����31��0 (c^�9X��d:$xN����9�l������ٶFF���TK��X�s)v�U�"���i��70S�+��8���Q�dy����*P8����Q� !D; �a6
�4�/ùc��2��ʰIU�Y����CQ9{� '����/��]k��]
����}1ms施c���R3bsQ9!�]�Kzm[�/Q�z��2O}��}��Eɾ�:0�ipT��E���Y�)�~���y��!��1��kU��]Lg`�g�cy���J�)q�HRf<��:)� ���x{E~~��S�:D'���[� `R����1�S-w"�фq�)�[��le�g��>��9
��ydSN�A*�0LA�H	ȜH�Ȱ�<LZu�ƌ6�l��S{��h�Ƞ�M�E�~�����y
&N/T�e�8������q�ko4Zp �8jԘW���p�#T���({��9�`��.}��d��S����k�<�I�@G�y�®��):�;��Ly��M�I�B���8ƨ�6@���_�lu��|�^�H�j-�%#�))mbz��LT�R�*PeFC��Z�ۥ��5��:��dwa �)و��z@3:k7��4hjOb#�H���m8G��:7��o��@zfk��f|�H	Oy,�2�W����9_�ؘ���F�}��
���B��2�<��P�O�5g�9a)�Q�	�@�gn�x�7�%Tf��e�܈L��G�3⫉E�&j6�1�YD�Ҝ>��B!ɣ�����k18&���aS]�@\X扴���0c[cL�zX�B	���n
O��^���#�8��ϴXD^j� ZpK��<j�@*����6�j#P4yk��{<\/��V��vRАU�qs�f�bş�Y +�R4r|�>��jm�R<4V<���j��M�iH<
r�Har�T�J�A:C��"Qy%) J���.����%�%}�֣5)��T��Q?d>�Va{��7%MbL�:o��<K�;��?~d-��zc��Z/9{#ΙZ��;�Sm�2���3@ep`٣�!R�7�%Uqbt��[�G���Ω�c��'U{Z�@�ewqq��Q� ���;C�`�,kn�Y-w=�$u$��E�ˊ��z=j��w���y��7}�|9��"/�֒5��g����.?����ТtBb#[�T�4M��qA���HB�acO	�	��ǃ�����CH�΍�T�ψ*N�0�Rbyu}Y�0�j�<�0�#�t�{!���m�|Zx���R��cq.E�
O����ߜ�ôpS�V�QB�v���_��� �W#���*d�\v�r�ko����40��o�k�EF���ν����:�,>�S�Oz�a��Q�0�b���C�B�)�5�L��Լ�$��їew.Q�qP	��ln	�gN��jF��H��@>zs ��)%R�OR a�my���?�����a�3W+�X'��~m�ȍ�Mx��š��� � \���^��!g¨4��6���`��^���2�S;|��͂#A�Lȕ�j�#n���4��_��������?���4u�;be31'�J��wE`�N8�aSJ��f��+����HEU[�(|���`:ӄf����$O}�ą
��!f����B�_��������xY{ӏ�̰��Rtw�4�2���y�_(ԗ~�w��x஼��HW0�ݯ/z؇��s�7���$ҹvN�@��^>�����B:NS����a%c�����R���Ը�@�ڙz#a�R��_^0�'��(�B��`婅	�ӴJ	�����L�M4u�@琩ڻ�l���$�Qy�,�HUV��x4�iӪm����0���0qx�K�)����<C�	�ܱ�3�NQk/$�VX[o(��N�Q��C!�Ir���lgkn�;�N��Щ�칢�M�e �cͿ�m쳸j�X�M���4��7�cؽ�m�j��]V\���lOZ�ggoT"o���*;�*�L�i�)�Z��� k���У(+�:L�+
�?�ཫ:�#�4�UH�!I?He�q�Q���bƁ�燚�ƙa(G���G�e@S�\�ܣa��' ��jN�����-�"��zʦ��(��?tމ�2mt�����9�%LF(w�}4�0����TJ�~�-;�Ih�z���A�R>�}j�L�G}�,��7��?�r쥨k��r��h�0�y7�����%��|R��#���kشH\-�s���%��n<:U�r%��oJݠ5��\�^�&Uݝ��LW(|I t�|��̤1w�9�<�at9�P�R���-�&�6���|qqi��m5�Ի���q���.���N�4~��bnP��\C��+�9˕?�}����2<�%���%����%���v�enD1���f�H�$�E����
{��P�,e FDn�poM'^Bb��vԩ%`�|T�x۵T����$�f��-�t� T#X��GO��ҷ�ٓ(i�yY���=�\)����F�X��%ͻ*��|�xt���6j����9e�g^<x�V�\��Bɩ�#AT�}5LGsd����a0��4��%�:��������S���r0���l�hF���p��yr%n�ԭf���$7�`�.ll�ύ��ցQo=/�<�m�8��d��dd�B2 wFͮ�A�B��L̈́>�|�=�x��Uv0ӟ�Hc��RS�x��1[Q�
 M'��xP�$5����m�a/�G.	C�vv~&���v1Q�g_lT�P7�;��2���Q�����TF���Z]~�j��e�����N'������������p�I�H��w�&`�-<+
�w���"�c$�I�����9���0���=�����/��1ڜS�*�Lo�H��}K�xx�����5O7��sԸH26;�5J^]��B�)��1Rp�kA�*"��J�7b���	�&>��</��R�z���s�'��ACjy�i[�����lx�f&й(4��Z:�GRn�ay�x�p�_�����tRϼƦLx@:�/�� ��#b8��&��������7���N|��'���T�,���(~�k��S��3;���bɣh��I��*%GoF�v�����3f��ǳ�3���J��S��£*~TkN�Eȉ�q��a�!#O���C�FK*g
ե�W�Fj֮�$��ǉ���bn����q�OH҈�����"'Zo��v����d��(���WY��S?�����h3�H�O��㚓Ӵ�q>���rE%���V>��& 6�zW�a����Ï���c��T���|���<Y,<5�&�ʓ��`��S�v��ԪiJ�]��#*}&o�+��,ғ�^C#�D�8�v���+#��N=����/�M˷۹],V4d�Ӻ����z���A����9�+�Ղ�5��}
 4��V��&��\7�c���ׅ?���4��7�'y[{[�S��c�)�=hܫц�XV�6x���H6um.�d���	�E�
�����7�1�A�,
6�$[w��=M�K��M5�38�Bg�yli�y�����B"��ڿ�f��1:o�1�<�B���%	��W��h�3EC�{:�K@3W��ݵ��G�˗%]�@�Elʒ���F�5or���õ�3��eBX7�Gl����%%�X�����9\�^@L	)�ĜqҴ�fm���TZT�t`#Nau��Z��=4^���v�FY�"�3��&���O���8b̜�ݨk�J�!*V�́_sٹtu r�G����1��S�vT����Y�#�1S��0�8�oP�#^]�R
�rS��~���`�"f����N`c����[�!��u��K�����n��PQ���!�����Vt��S�3))|�k�R�P� ��d�q`����P�252���_����y��2� 6$�ᙑw�sC�0�4����?���>y��
�b:�f$	=	�@��8Ro�I��+R�s볽��я�4�N}1����*%�*J(���o�����t������67��!2��Q�X+�2����g(c��7�w�g���rS�	1F�G�S���0'���xJӧ@�]�߄�wW�W�P�G�Z7:��Q��E�: QfB��[�I"zS���065�8/2�QZ�1��u��԰����=*�7*ލ9���Z��i�,�Q�c��U��P��h�7 ��zMH���H���{�&O�c,�ʢ��'	��1j$d��!u>�f|��50�ㅃ���zOX��S��/�t�4�H�a�ǚ4����*)<���@��9�U$�0������y`�W��Fg�6��nPk׹�.p2v��oT4�	��%��u(O)�|�Nuը~J��wV��ꃈFI��,OW�bo3���8.q`���s�u����yσ��[7)���9�)�j| �4�1��7�,o�@�yI�[H�p�]��9�lԮt�� ��z)�K!�Q_�Wm�"(��u�߰��@��#)�� ��8|E��+='�ֹ�q�*#�Yx�����l5M��xz2�Ϯ�+;��S������iB��ZRka~kʁ%����uf��y0���K;VBy��b�}���{Q�ɦ��@�'[���rx㚜H;��%�F|��C�3%M�
Dw�a�3�rR�x��]gT�Y���QG��X���}'2"Q������,�m�{)'?��l�V����T��H����Fe�@��B���j��q~z�9H�G�� �:���J'U�Z3Hb��B�R%�υ�A�TVd KO4�H��d͆CE�:{>-͚��2�>�Q}��������b����@@j��f<{�9��n��9i�M�Rt����3����i;Vh��F�A��b���q:��#�I�̣��%�16:g#���!���#4�Ws���V�/PD%
<�����|�b�l
�43J���B/P�MM���� @�-�:H��D�L�pd/�ʫ��C{2eM?�:��s�d��$W�P$^� ��.U-	�̶��I�Zݟ/��e�r�Eǹ㾩J�X r���g	��z!�	</*	0�닺��i������w�r�~n����.�xGO�	M}n�IYB\W��>-o"�ȸ��d�	Xڏ��Q�C<%��Vx48�8�������.��6�H�^ƣ*�s;��Խ��F�ן��>Ҙ)�Ϭ�tZ8��_;����Kܖe����a�Vc���X��
䅸�=j���І(^�7�q㺬�$1禇��g;ο�t���[۱� ��<�xq�s ���%�Oy��
SΣ�!ՃeO�0V{]���X��$������{�T>���Y�� �ph1�k�zT�C�*�8p�c>���YƲ�;'׻J��jLΆ&B���7"��Gw��w��r"ul�Ԇ��vkt��� ��M��DB��1:o㧄�����S���r� ���D;u�o���D��&4י�4�S��F!L�	#:�j�~M��#�J��m���F暎�77�t�E?��!���iI��!�RE9Ԏ����e�ݳ���96�2lp"gn�`{z�lR�W:�-���6V�l��Ƒ|�W`I"bШD1���^"j6��ֶ��u��8_���(W�I-�lV�^���%Ngs:.�AYq�ꓛK~ u�)�.�v�ۈp�x=��v�YnA�GrQ\��H.��1�%�y���w��(�8(��D��D�ɑI�0!��:#Ob��w��<��X���-�`�� ��F�N<{ri��X0o�&��F(��)6;��py����o��d.W�4 �a%��W�h�w��T��
a�B�#�.F4 �֒�k����Ӏp��\�=��Vn��� ���1R�=	?����'Ԣ#3A�5�4x��$�gs�zj�7���`��쯒� '��qO�mO���ѕ�g!�vD`s�
���r�P76
��58(0|D�\�Fw�JىSF/���!��B�p�;��"�,��u�h3m�I,E�WNv+dn�Áq���J�0�0Zl�*��u�q�s�)�Χ�c
63h⨀�F�3��^:%V�6�y昘����(��?�8y��uvvnܷ��:W;�e4�Y�۩��\�޿q}�fo���\j=,���%1��Wo#'�!��OI團3���Ta��z%C���(G�	*��Q��<�+R�
���6;�-�਍H���b���&z0��r1�)�G�����8�"��p���{��(��������ؐzi�*A�c�G��9��ƥ?��0�����;�����Ճ�Ҁ*jSM�<�u���#*Ž҃��b�%�<p(\�$����8".3����з���������Sz�~�\1��k�dG^�t%MQ����z2�f��!�oDL�*�� ,������꩓��%ϳ�/�3���Kt3�8�籔��}���UT�6�#�I�C����zg�
��m��!5Z9i�Bq��j�g�ռz� L�N��˅��~�*�lfׯ߰��-R���<_᝱@�p!�S.��(
��ͩ\�u���Q�F�S��U��gmB���5����&;�uԗ�x�ao��[�-�?q{�	�V��8�JTJkԏ�"�6��^Fe%`�Um��ޥm�ˉVs\��@�ER�YSŊM|B����1F�Q2�䕢R����//}�f�}��#�:y�TK�E�������9)@R2�D:�j�/ۙ��Jڮ
e*ok
V��ig`\��[���j�1���޵G�$���{DdVu�����Ka�IA߅��`!,��Q�R$��=�U��f&?�k�YC�`f��2�nv��s�9���U���ƶ��|{}e0��R�K���i�yPR�܎-�������C�`'�� ����3�ԉ1�6�5�����t�L #%���Տ1,%�� ��#C��L��q�ʕw�ޟ�9(�*�6 f�ո��7��q���s��R%�+�?��v,�Xx}�^=�u�;4K��n�x- A<ቴ�������f��dK�D��%em>Vt��6mr��&�MC�~�ۅ�,�렐�ۋ���%:Q��W��E�Bi!W���
/wH 'ǫG'�i�s�,�[���&k5��Oϳ؃bmv�v�k6�;*	m�!V�*еk&��a�B�����Y��'Wy�2�� c[��(s�n�N����q�@�QpSk���H�#U��z�#�b�N��Ƴŵ�㡃$| �,@�w��~�3SzF�s�|&��Cw~G-��L�z�Y
��﯁����5H	��7�i�U�l'���xa2��� 2�~��qzG�~�s�k�epm�?r���A8ݧl� �n|ʮ�\�z��r#�@�,���ܙ{7�a��r�<#�e��9��37A�$~9s����;����J^���������.X��&��Wd/7.�Z����ap��p�Iݚ�쁡��FiJ�.49H��v�p�l7g�M
b��/R�9*�^�|�e�ӊ������[� a�x���.s����+����!ha���W9DCdB�1~�2�Ԧ{���O�����<��7O��#jO�+jeA�� \5H ���_]���<���D.��٧#�,n��ں2�ŎK5� ��LA��(a.Qk;Μ����߀
��X�ȍ1|���ݸ	�Y��u��e� E��L�,�J& �Lf�{����<��e�J-l��>�Z����0��YKΡ/AJ�(]�2�A��?'�Y2ooֽO�Gw�r���o<h��Ip"|g�aS��*a�=fe�4L��za���HO�.
����֦����	&9xF������2H+#��~�zO?��S�MJ�����v	�I&�M�T�S_�~q�0]��}Wm���E�!�����ӌE3ޑJ��tx�%k1ז�¤��V˲��`���~��5�5��F�UXǴd��kfa��!�.,�(���g/?��ʲ���B�">�u?I�r���@���}*���A�V"��w4�������&GE-9�����kn����i@�u_��J�~�k���4���,���帆�,.ks�z1��}�]��X�5��J_�]O���pj}J����n�E*<J�G���-�&.�E�}\�AD2����DI�kl{`�j�<�]�c�F�h�&�5�1�-� �Xe-��i�D�V�Vo�L_iG�g�4�P�BU�֬��D���}�]P���D��Q�C�&IYe>��B)<�(�jʨp�����hߋ���!|@�����������Cqz��NhֵRD��ܰ�Cm�y��i��T�]J����tuQԒbZ��p���I]�ԭ�/ds����37���C��(�{��r��\䂺��ă� ~�o��gs�,E`�$ox��Zn`�����[�'Eq ֠܂���LU7���y<Q7����gvZp�\��}�1}\O�R�I9	t|��\<�$A�e��17��"���:�,��M砜����}�?FBX@ы]���P+��M��s[�"=��d�Z>�m���LmL�0�r�A��.�F���@0T�%i]�ڕt�����M�u���˓��]����Ey�*'о�6e�#I$�������-�9�b�^.⮌�M�RX/L��א����,���9Hj��N�l���SܦMփ�6������Ðu�,��~hK�A{��	{T��+�r���^f@X���]���w�4"u�����fvj(k�:�|��8&�Yx3���F�'�һpN
Z���-\�23�N"; ؂�#�{�^9ve�̜-��JR]�L��z�*Hl�7cr�y��&���D'���S�H)p�ƢA&��)#HcHc�gT$kDp��������U4p��dȊ���:��(�8����[��<Q ���1�-1,��plCW�x�7��k�9Cu�:�0Ff��Z�G�e	Ҳ5عpo��^�\�_�rtg�u�J�C^���,��U����Kz�ǋ1�͘��H������͜�;JZ=>{���ϟ���֝��$��E�^o���&([N�;��m2� :�ڎ`���On�0�SX��f��@W�����^��u5���!>�0=z�IY��æÉ �M"�@�qr3�~��_�ƅ�����u0�T����h���ڌ$���h1Y}7��ϸS<w3Xz�����#�U�����vW�c���d䚛Ph~Y�3�g���t���,a-3_�X�5A�����l�M�v��ybI�H0
�� ��NdAw*!����"d�t!���'aV�I�Ǚ�B�����7�_jK͌�G�5 �PM�n�I��7k|ؐ�r0�\���8^d�`�e�ȑ)iO�-�8��fkO70:gL��OQ�z�}��Ί����b�'Ye�(�斟�Cu*��rdܰ��讴�I��Â���_�|��-HSOdn�0$Zb����}�\�-H��Gg�z���^ �|�(s�e���1й���&+B�l
�*]�:D�>��%3͝5 ��@~�����Yg�X��`bR���J%�?��?���>-%Z~�f֏��C�U-RB��襚"e�v�^HRJ���)��m�i	�Z��D�Ӕx1&~�n�Zw0��3��pr�^�."9�I�?����T����v��=�T�4�+HVsx*��H
ʡ�d���-�l���,�&Ga⑨������@D�^.d3���,& ^�j�&��mZ��}��">�Ki��g���E̣�<�i��e;�)�x�yr1 5�ƫ������^n|X��/�	@�g!���t��E�S
���Q���U�[d�O��Cf �蓶�˚�ʑI22,>�Llyrrl���u��f@\���T�O��(�W����Tu�N �?��#�K��UeF̪��x1];Rea#(�Q{�7Tcڹ�}/6u�p��#���R2�j��9K�A�A��Hj��Q��,w�}�~��~����?�{���E�>�A����Rdflۿ�g��4��'�w��g$j��hA�H5I��K�d��N�=��P���y-o��� nh�IbeW�(� ]�	����i�Z��V�qt
��0A�ٍ�#��<�$sO�b1d�[<J�	CS��/z��V`̒�ږ�A&Lx��	���y1��#ߚK+�;ى�
9@�������JS0�4�G��"��@"������E8]���g��u(�J��AKn�{l���Y��XMAi������~�8���yY�-6y��7�)ň�h�5O[{�|Gބ�:�>M,��\�PH�{����0h@�����!�:b�A��;IKQ\Z���:���C���E[V]'&�s�M<��u�l_=�=y�Յ��K>� �'�k"c���CL�c��������.��k6F����7ls&��z���Oك|��e��0�,Ԃ$�p����ps���g�7����0u�Cmp�E�9mͼ��+�a*k0�e ?���0�?�����Xx���g�̘?�9>`٭�BC������D�r����P��5��J��ًG��o��-b�6�uˮu][w=h;���#l�T]�Ј'��đ�8X�%�s�N�-�/PG&u8���1k#Q�@�����1&1�$���$?�ΓMl?���ǻ@a�؀{���!!�RJ��+;L}�|9�6�!iH"�]?��1AP{���^������fU�Ord�m��'W�im##�!v�\G�j)�ǁ@��Bք��p)9���[��Ռ��0jn��󴔠�{=���u����̗%�y��T��d����vI۾�@�����J���qi����)6��V	��۞F�p%gkáTy�Ae�m\�,M4�G��FFn��l�M��E�-�(�qˈ�ȋG�����țH���N-�A��Y�=lq��j8=��B*,/�b�uQ�'y||߂��:# j-��,ǝV���Ό��8�����Cv��P-\���� "ت�HY���l�,��g���\��$#`�SYL@��� ��
�(+��S%Lޚ5"]]�r��<ɓ��M�1�۴��4����U�1�^͸�����⽊�5(g�Yqku��	U�#��G'�j��,=s|�ݟ�ﴺs�@�1`:��-���!�����pW�1�h�Y���X̲0z�"�]�.]W�IV�ݢF:�� ����M8	�������b5����n����޿���?����ٞ�d�.�8�r/J��W1�u�3'�v�O��������f/��S��'$�2J��h�<���bb��jAy/���<���ZL9��"�2ܔ���!c`��u��z���=�m�#IFk]��:�ٹ��z�E�y��� �y��>�.#�.Y�ze�3 4�)B�1	����S��eۦ�(�8,̴p�y6C�b���1]��F�d/�>ݨ���$g�>6��@�J�L�Ɓ#*�M����nك��U��ŸN��t$/*/P�`�ca�P����h>��NϫL�FxP���M�`�m����~?�%�F�~���n�%uYD�B9z����������ӑ9%Y�ѐhL\b::��L��wr=�coq �������Y�䲌4�ّ�&�'Ax�r�x��$�|��4�& �0�[��_~I���}�����9=F��-���Y�3Ol���\�حkô�u���ě#��6A���6O���&�ԡ|������.Z��k)��fE]|�E�!��o�죻|H�*������f�*��1�KC��N%�]�?}�'�ʋ�H0-���7@�`Rь��b�>��'�.��W�@�h�	ʆ^���a�-�=�:l$��`�Q$c�i6&����,�3v������4L��	&��ˍ�لA]Z�m�K��p8���|򻭷8���l4�QPA��=Rk�L`���0��R�A3�"q�!�ޯ�u]۳��MSTf��Cɓ�sW�@�Q�ib:��b�	K���W����M���<#����`��`&�e
#	����l�Ę��_����fv��.��h1��A�c���	�rK�u�����|�b�)��5y�ˌ<L�aT|0z!�G�~2��L�Fp��]��{���M�e��)F�їٳg�)T��S�J�W�G�h5�&w,ԃo�L�;`�<�}��E��*m�R���<��hU)�{�w�u]l2"��"i::�2/�W�f�Y�=�IJ"qj�v?���A�ÍTfz���=�=I��X��)`�$LvY�kH��t(NӁ���:iU�5�-:����`���|�+�xT�n"��:?k	�sR��$=��	)*3�V��B�yݳ2N�	���B�UV�x��r4S��F@�B��������	k@�鍠��=��0�%L�Hp�2l{��[�j��$|N��(���p�ڴ�#n�0�9��{��2�)�}� Z7���9�]��;����� ��~J����i�ݛ�z��!6K�����J�n��N*���Kz���[�`.|�����{��"���v���M�'Ϥ��IK������#���	��ì�`�\:}JN�?0��B}A�,�r��ѡ0�� �<(O���/ڌѶ���U}Y�]�J4�7a?ƾe���z��&ɰ��HjO��+?�����aT
65�ԷWICѐ/7
,�>� mАe��&�	�D �b��ؠ{���3^K��ۃ!�qr��59l��Ǧ ��m����p#Q�Jҽ�xx0��9Z�������kb��o�]�.�6��W�*��Ў�9Ԗ�ƪ0�ag��S��(&t(1���/�0��i���w����A�b΁,Cm�$�x>aswt�ݍ?e��q��d�r�}@o�!`��F����������H_�_xֽvD�YJK68&��4%���rd���h((�����9��F3Ȥ��=�|$�*�{ݟ?�5a/�P���F��C�������*�s��l�H�h�����B��"�q�$�l��ωړa���y�h�*����bX������	(�B�r���Wg��85[Y�����̍F7���3c���7#^�d;���a>ɓœ2�.��4"�b�t�)�#��R��e�S,$�O�=��~�z��2��J�a�+��J��LД�� � C�
�ɲL>���Li�e;������ϟ?3�)�t+�+3��hP��[��v�p��`�_V9i�B'C2�'O����6b��h�ـ2�=GF=�	��XyY�7��c>�J6'�6(PNq���������B3XXn�P��Z�|
�t�a���ߧ��~�D�a���������F���eO�tz<5�ݐ��C��V�߀�@�B��qw:�������\����/��"�X6�9,�#p�	��㏂ݷ����b����>�ͩ���0���!5�������J~����(�8�M�j�$$��c��K���(|��>�P�1��[ң}����z!���q&$lW�������I|Mrc:��ͨ4�҄��<{�E�Cɹ���(9�S(� �h��:��]�]fTR��׬���l��(s�!S&P��?a�pr?I?��N��g���`����i�6��~��n�W�P�� �����AJO3�_ØJ_�����m���}�._�b8��/v��j��Jp�g�x����D}���l��h��}��V��y-jx��!���I/�i.e�/�t��:�o��Y�}��/�lqb��tvy�
8]ג~����)���;��n�Pe��z�Q����#����8�.a�yl.n����alw����#.:8�!c��v����Y�����(ҟ�̱�#|D��-,�[kS�;SX��&Ќʏ��D���Ys;%2� ��}���:��P�-7���O3��D[��|�$�s��Xfք�$�3{\@�w@M�iě���������� ,�y/'}l��pc:�܍H��hK��kMG�����l�<��B�T~6y7[��>導�?�	lh {����MA^��p�q�"��}�o��
��ӾNf̠{,��t�.�V#p՛Ā>1����	y)�'6� |�iz�fn�S��\S���x��!?"��a�H>�?�.�J3�CS��P�h�6/����1����ӿ�����(�4�����U����?�Q�W�'�y�r3�߭4WJ� �����2��,�@��4���Q~�	���@���<�7i�����T6)Ӄ��H]����1��l����a�X���c��6�HJ�R���k�R�*s��ܓM�b>����'�u.��4��g)�L��0��
���ۅ)�G���YX "e��t��pwN��8��>�D�y�T,=�]�J+�'l��R&\e��M��e�m)D��n�����n��������F39�ईf��El����"b+ �!�i��� �0�!�C�j
���`3*�!/��ܳ��A�%��r��M��;3$�H��F�~�&��ۿ]i)ضR�I-*ң�ݗEL	�&R�
���LhQ��Ƀ�a�D�.��R8�0v�ߗ��� wŃf�'�t0���S�s'��Az�J"���?q�
r��N��.UO&6 e�/�y����Rk�o��?�,�X,%J ;<�����`�ˌ�.cQu!�\��q7#5���]jѠX���P�H���/��ߘS@F��)=�p�<��/�t�(������̓M�J��'��ۘ��:����}{��O��Z�[�ow�8��E ����$H�{/��k�V3Y�n�c�	\�~�c����'e���^'�]�Md����]�˾^�>�5I;.(�%y��S��*���$��#/S��C��/A�j>�\r���l�yװ8T�'SS-Q!QYu� Z,�������~���^�1�܊����������l����4�nЅ�������e�"T���&~��L�)4�6kNa)�`| <ͅY��v������w���<#y���x����;���b�Yߑ������V���8������I)����͉�ɥ��@�pITn�G֥)D��������	�9%�k�;3�)����_F'��-d�ϫʼp1�����=���ub�Z�D*;i��u�\����/t6Zl^%O|X�S����NQ�a��EY�\ZP�`('�\�] ��$�9[�K�������O�i��=�b�7U�s�;�L\�7vgP�8/��6�"��R�s��%J�A{���Yte��b�m�l����sRh��ϡ{U�����M�M��f��L� 3=Q#Z_	l|�j��J��NLI��<�)�"��ҋ�Ϟ:K�!���7ݽ{��,�3� ���N�A�װ�*p��a�6�RQ�1���1}�d�?���j�(��߭�L GvӻO�'٭�s��/��z�����,�}r��y��-)�����������+�xR7
m�J]��n�#Y?�I��N^�A�H��L�9�gΕ�In�lވG��v"�c�)�����(gy�v���BXO�!��~:~=�H�ݹ̌oN X���@��46��/���$^��A��qH����z�|��Ĕ�̭���22���@i�3�JI3hӢ`.���HhK�33@y�ރN�� S��,3�C������PͶ�٢�>���EC_�������o���?�~�k���t��N������Y�&d�uWЏ���7/~0�M���@�bMڣ�������B��f��9�6�ꦾ�������&N3i��P���Ϛs5���R%Mn LX\���=۩c�&`�M�q"�!t��ܞծc�k���	huW�^	�w@�W�a����Y��Htx�Ц_oWg	C��"�Jϲ��j6�����eQ�e[��L�N�n�7`�89�F��a1]�|�c#��-��b1�0x&����XY��%�Ap޵SbwW�ﲟ/�K���u%��Ů��]�����)
�!�FZ�����-YB�`I���Ň��Һ���hB�4P��Iĝ�w�D��AU�jÚ*[ǅ��4&RВ������+��u�H+?������k�2��A�&�`l��+ 7#܆Fe㘲s}�B:.Z����d�P�~��1}9;�Ќ�Ren3����t��s'�|16��%����x})'�HI�R�����	ˮBa��7�S�yO�Ncݣ ڬ� �=��ނo�ɮ�5J�`�%3AQN�\\�M5�s���Z���@t�9��`��(?C,1m��ڙ��r��Z���°@*"����:�i3E�����3�L�0DH��\T"'�p�r?���q^��̪��\�Ϝ��"��:yo ����=�/�y>z?�"}0.�Jd��'�1]�hJ�u^Ox@�l��X���U0w��ɒ:,̌q��uM�˨�QM_��Y��`�.�r����9�����Vҟ��o��C��c�=�I��ʗ&�)����@�c�3�x=n����&�D�v�K+���OM�`͔�Sǳ�QN�z��������(�]�˕1:�荇�c�XPhu{3�N�h�/�����J//=1�22-�*iB�-��-��G �I�Għ��4zWz�!�~R�#3�����`����sq�I;�)��6�X	 �۞I��R��h0Y�Vz�l��F[d���͕C��Y��/�Qfx�-���NkIX ��r��O)��V�s�o_`����$X�	�{B`SCm��,�\.fi�J��(�~����j��17=�B��߿�"���Pǘ�=��7z�)(��n��G{t�P$��H��!I�fI=��7���n�+K�Ȋ�qX�9���y{�*?k�rr�YgG�&N�aZ��>�Z�^-a^���c�k�Q�{�Q}ůc"L?܏�(�d�6%d�ɡ�g��(��2��![Mq�m���?3�NM�T}����vP�`�75�����)"S��!�B�5�Wg�H����]J���xKl�pvi�k���$o��`8v=��'��`9~��V6n��dԊrܒ�p1f$Iuw >�E ��${
ۙ�ؐ��j���\�hsDG*�����r�|Ն�xĲ�7�XQN�Y�~�Qr����67Cw��g2-�w)IsvV��%t5צ��e�_�	��<l���A=����s}��.������������'�;�+ŸUO���8}�l&0ۡG{���<��h��d�W�t:����x-��:?W���10h��e-��g��`��s�����N�I��Y��s� �_�������Ǔ��4S��X��<�qeQt��7[$-�?M�8�����7u��[�4/�:Z�E�9{ʙ�Ex٫���E7���=�?!;���D͉ڴ����5�˜ �@��E��7����w\$��Җ�7u�0�j��" �#���\�xr��=�$�yc �,�ҙ�"�#���q�ʼ����"��`��8Ъx&{Lr&�aQ8lU�u�4�̢.p���FЦ����U÷؜��G����3�ڢ���b��{��x��:�m�]�瓙�M�3�9<'z����p��J,o��4��ݑ\�Yx����kwV]����c��wf��#3��ղ2�C����6rO��k�LL�m�3� ��Cf2w�i�y�-.ټ�/_�p!8���$)Fŉ�f��禅�d�67�3�?�4uߘl�=�黸�#�`�	M�k��7	�~���p��z�s8���{��őyC��P�E�N��M�%$���B&�`�4�o���^W{`�%�m̀��k`A�ɇ�ve���nQ_#�ܐ��n�f&Ǣx&�-����2p�*�E�|t�5{%%|�q��j��Xa���4��#7�M�����O%͙�.���M8F
`����N�Ӈ�yV����o2<'����m��a�=�[���=���xI].��J��T����,��+���3��	��A��T�Á�=55�k10��w���v���.���K�Y���Ad��1�)d�//) �(��x�˷[5ԮA�R�w(j�_����7�Q֘��c��&�('��)J�m��yF�������g~6���ӓ��Jװxn��nR���< �wZ̺��Ԓ��
Z�N+c�=�̛�����Q�>�΋���a�����6�\4��%��mF�Bv��Y��t
��F���)��܏ҧ؆���H�0�%����ẆΒ`��m�gS�F5�t��Y���J#�� |��5}(�|�v�v�Ȧo�`��Hق>MrC����gp��eyn���tF
\�Ja�v�p)l�Q��g�g�Փ�䒳Ob\٥D���q���J���}j��c����(#f�GE��h�A�sSN�:�X��f�!M��X)xT��$�Qz7�5lݙѢ�K�5�5�ck"g�s��;=��#wɧ�K�O/i��fvim�nh���E��ؼx��w04#�}d���Up��I��C�i�Պ���fP~���lO�����ex�sxO	`�S��o&��@�4���݋2�����d-њ�"��z}���EI�Em`}�#JW?�w�T�uއ#x����z��)��i��y�f-ŉ��AW��$������ͺ�C&����4;tv�_�A5�Ѥ*�d�ɩ���}�	�UЩ�h)�qS�K�{�L4�x��'87�W��q`��#䚅w�BC�_��#:��AB�V'�3�l���M��ɜ�J�"XCV�'��h���J+Vk3�#Z��Q̈́6>�X�
2a��-�I��
6������>T���8��"��Ų�D��h�䯿��F �o��oӿ���F�$����0���f��b��I3 u�yjr�qa�v`j:�hSv��h� 8d�0��liJ\�k�v�<��K>աI���Q��)��!�|��F>|U2��!�Y>�� ��t�9��[#9L���%�O 2JJ�Ҫ��ʝ�ч�Z�VU�����pq�s#�����ɚ�J��]��0!�@�7F��z���dTj=BX7D��w���-):a/X�E#KO���ɨ뫀5��p.+�`��z�c#SqN�8:QYd��*T�x.��Q`6�*��-�9h�NtD;��o�;S�L�xԡ�g��p'	
XV�(�>���v��ڦ5I���dJ������Pch(�;Gq��;��J�ǝ��E�X�5��X�5���f�A�J��>��,�<	�}�.��G��HO�����2 	���wi�%V�-��� #�\	}H��)���:�����ڭi� {�-�>��EbC���hC��L�,�P�s"Q�w���@����1{|]�S8�ؒ��\����'_sYг��Q�b�a���Ua��̌<Yב�~}s�qQ0���k�Ϲ{�}xn`��a�n��;��S�W�70xl:�էH�9�/�ڣ�a����
bP-.u1=jxCy�
n� H:�8	� ��T�Hy��x��c�o��/bo;�Fi�Iߍ��}�h�'O걱|��d."U3NOH{:Ha}2Z���b�	�*�^/���҃���mU:�/�w������3hc�HL��ڟٹA�sg0�F���Fb, g�pd�k蒥r�L��H��eC��Dj��{���o�����5M�R��GOP�-�
�mLa������]<�D�8��F���"���]l�K}a
K!�H3@���Zې�x�'�O2n������gn�_�5a��T�Tƃ���Ɖӎ�I�}1��A����}�	���}�j�]//���ݜRȅ�]��Ri,v^��(v�UWCS��p�5	E$�mܴ~I��w�$��-`F��b��ً�����5����۝Ư\z�d1[ �P�Z�˯��lZ�J/X�6�,��K�^�e�IL�p���/�nL��SYa~�3(궥w�n��cn�`�b��A0�ڞ��0@B�F������f�6q��>�����%=�捖��F�?�@�w�6N�϶���.������$��OT��D_\��9��s2� o��`�ll�%�V�X���z >�2b��3>�U�t��KJkX�ؖ䵩����{K�}-Frd���l&�D��F0� i�=�PǗ5��"U�'B�Y�&AS?:!,\57 q���k��0e-f��4�"K��=�)�2�����񢹞|�w?�"o�k���j���ߋ)��)��d��!b[�3or��")���!ƢaǤb��������ě�� ��56c���ݺfc.�T��-G�A�z�i�C��]
 S���IB���KRn��)Nn9Z��6qP�u)��.ջ�n� C�b��@���kf#��q�����R�?�T���F*&_/�߷x�7�" �ي�	�&/��I�B0Ƚ�.Ob��]V����y�ﻯ�G���Ej�:��zYo��q��Gef~��T�M(�l��4�'���=�O��I,����5MN��Icrv�K��D��Ez}��ԫ���[�ʚ?kz�����QT��ӂ�P W��{� SY���̾���&��%��ȸ�/x5�"�E�y��Oiu����m�H�̦��+�$N��^r �<w�sS�����玍��lU� j���t�`��{�^8sK
5�:C'd+��޸�r[�`{�23+o��ŭE��EPmޕ�v�����䶬͆���0�їv�lU�ٔ����|O�N�'����]���f��k1�:�Q�~M����������.�Tsf���/�]tP�r����:�3���7��Xс�{��"����YЩ_�)H3ۊ֡��춯�+aio�H ��K04!NaF~��i	�GV���8�u}���.0a��o�A &�&�%�=�	���1�\��P��L?����7�!O��kku�w�zSc�#f�@܄�q�C6e����N��7�bu�~�aH������.o�T|i���2)�(���M�2�o��i��'֙�듭�*5�����c�s�?d�8��W�v�X���x|[�T�iQrs�_�p덾0P&��.��en�g@&�U��k�/�q.D����-�>yi��x^�=���R'`:��=j>s���EȊ{��"^��w���\ebD��T �v%K{�#�����1�mhj�Rx�M]����N�-4w�C%j)㰡�)2["�s��|n(է��ZLW\.qW<�Ǹ��VtU�ۏ�-D;Wmj�ޥ�Kv����H�>e��~$g�I��t�t�� @�@l�e�����L?��ڰ��pm�'C� )�$"~-8���OHqxK�K�t��t4A[��QW�V��T�I�Xm�Ɠ�]N�c����V�go-�w�ky���:�.��W���o,Pr]9�Q<�~��Y,
(�ͦ���lG'��\�(4���q-)Ͳ�5{�~����_���
�2U-М4�v�j$9��4���S�$�b�n��ȆJ
{�ɇ  ����V�3�X��~��]d!���fm	�����)�	q�R������.�Z����Ǜ��U�d�I�DF��ZE�z0��gx�汥���q�����j�a�Zm��� A�vU�o�z���m���%+b���V�8��Ю�|�Bh��/D+�����o�?¬x�?��T�%������bӂV/3b<��<N&��(�o��������Z�Z��u�=�}����o��PnMs1��:@6�l#7��t��	(؁��4U�O���3�w��9ە�~5; ���8o���x��_Yܛ�B�CX�-E{q�t��֫؍#&��I C�	6'��^��c�I�v]��&�3SR�P��G�����Y��9
0�gIj�-9�a+��*mT��Lf�T<��Dv�3'2�<�UF�����}�0�0�U���:}����}JS��wr��!2V��)~rP&�|.���uyJ�5�,����)��������tг�Ңs嬯S��%���6񪌢7u�:&���H)|���86>J�9( h���>23�bpХr���l�=� ���{2�MA�Y�}<�.l�H����,W$��̚n�:�	�=@<4��ڀ%�b6[g9��%3���}Ii���u��GV���#�J{�
<�a3<��ݎ��ޅ'N�P��~��Lq���w:lg�C4��B/��wM�ɸ�R� ���P�,���?�ʹ�$�M����`�4�����Ugmנ��y"�Y��#�.}�]�';����`i��4���߿�M-��Q,�D�5	IG`���{��&T#D����:��c�m�(Yx�ų4�Z8!̝�I�R�dՌ�R�b�`�q�������%���ٰL���M����6d9�y/��XF�1�A~9d�s~�i�A�/hK2�}��eʷ؟2�q��� ������/<�P�-��8��n5���V������l���,^`qH�&R�?��>�+!�8�pG��/e	�J(��8de�ؗv1+.	�(�V�R�p�R7�ިW��B��yr�;a�Y�6"��/G���i�E�S]�d��8Y��pi'dz�2'40![� 0�m�̦��v����ፀ#p�8z�T�u ��\��Sd5��l~�����i�]�0���U�jY9ُk*�	��[�N�h���v�;(G�Lɋ�L�N��k@�)6ށ��" ��T�o1e�DJ��/�4�r#�е٘-�ɞ
�W�����bA��}L�Ee���L� 㶲C糢�i�D��U��R���>訜�χB�'�w8�ꠞg����
Q�B�'�4z~.YXÓ#<]�X����,Jl��՝Ё��,ӓ���_�hn�M�W�ڞ��`f�̔�6���� E�<����"��������������7�ږ�V��ḥ5ե<�[n���p�1ka���ы_��q��]W��O!������M3����br��i���4��"���g�g�����|��%}��p���9�k)I����Ґ�Z��=�qs�Whjgh�{(��4�ӛ`��2e&O���I�ݶ���Cӷ�2ÁJG�,`vؕL~2�#h�K6Q.�#�ބ"�O�����0x��^,��gA���M���6|%r
B�躇�6u�x��f��}��E��I�K�7$:5�C�.�t���nƅ�;�pJ��1��JSȔ���"�5��|� �A�O���������i���UB���]w��/F Ղ��I�(�W������bȊ��lI`�u��bccSȍ	"�r��{)����U�(p��#2Z��I������� c_/�Á޾>ٲ_��ۚ�����O���{,������?�4A=W�I�i��y:Pzi�q�)�&g����>.~�p}�8�*)�X5����q�#���<�e�5O��f��5u��y�Oȫi��'f�:'�B~=D��T���f^R�<�8�$@J���@B�H������_H�-��kML��Y@'��~�p�a������5a�Kk_ɀŤv*����!�tx��1%�
^�}2�����x&�ơNP:?$�F<�G�N�`a�����6µ���C��2�|��vN�� �~�i��<�،���N@z��� �C⛷��7�$�.��2ߏ������⮛�M��߿�õ�YA��~.t^���D.jO�KY���� �.�K�+ۼ6q�����BY���������F�SZ���=AN&s(3eK���7��0��?��um,j	xr�)�%��� �����1� ��Lq����n�H"#(��??�8=LT�F
V��HlS#b���Nf�a��ix�YY�[q�g��^���rR:���VJQ)����Mm�$��=�3M�"�9�:�J�C'+�<����H�=MN�ExeU�N0+u?�q��:u��o�ȶM�ѥzzlv�҆�]�B��>I
W$��T��K5�J�C����UC����I���0m������Ǒ�.JQ����,�A���>9:i���Lw+X����,����b���4a���Øu�6N7+v�P���H���q~4���ܸ�@��4�ȷ	�W�����;�H?�� S��  %G��o�#����urSMT�dn�+��.4��3zR�ӷ,����YF�'Gg O�g0Y�^j�DP}^��F�?��ߠ�\��4��8�koN��v7c:��>?;��D��	4Α�S��g:#ۇ�>�^
7�{��p5�s��ƥ��M�mi�8�,�M�#�~��P�o�M�����,��'{������'j�����6�(�q���[����%&���˜�fX�e����J%uv�W'0�����m������8-�1` [�g��}�a�1�0J���3��]*P� ���@�>3A����ϧ�D�y�idƜJ�O��z�#�{2�vk�7��(X�Ӑ�����Z�s�m�N�c�lƇ�ʊb�^浑U@�}�=r����e�?�����]]�1��4dn�<��2���ȍ�̪�nu�V����=ǭR �v��\IރF&ŝ��N)�R/�z%��U�+'>N�$`1�tGתJ+`��z�M�K)�z.(w\?�]d�
�H��굞]'���e_zj��`ں���1���@�%~�Öt|�O�׫i�!<��پ0wo{/��Fu̅��x��w`=�L���+kA��l�,�W��Ee�Z����ƽGp8���,�G���|?Ƞ	ٺ'����g��s�j�>��<x;
�0$�g &�v�c@���l���b�nh��?L#ה,	��R!����#�=5�*��I2�c�07>�Zf�4[�I؇���-������ɿ*��Z�5�4�o�	&��eM��o���d^��tt��,�����l˥ �X���g��	5��cl[Ub���Fj�L"��Jst �OP�U��l	:�8�ޘ�� ��H��u�ѹ9�%6Xa��t%�M����������6���%�Y=���g�
���8my`�Ƀ��� ]���tٲ���Y\%��	V���
��])'J��v�qW��e֛'@��S��cn��'�\3�Z6����T��i6���md=K��pN�I�{�K�����F�#l��,�BR�Cv�=,��S��nq&ZVo�Y�[�s��p{W%������)��6�ʆtMĬ%��.3ma�G8E��>�����R�j�r���۹�����<���%�}+�?@�+?�1��a8Iٍ�u%�'q��"��F/��~r�ǿ����z!��ө����w�8P����t�7�(Ĕni��	RfINE�>��ک����y��Z�I���^�YT
~V�p�MM��fEDbA��M`P|�`�������q9��{ʅr��@��P�PF(�/]���[��~�Vj̕����t�d����p�s�.�U+Y�Vj�Έ`ƺ�g�T3#��9��fѵEV���L��ט��܇%��c*襹��d��!�f�qsn�l=����-1*@���p1����k�G�MX �	Թ��&���F���M8lǝ��Ff�Rg{�sZz{���2g��~����%�֗ݜ�?��E�3I�b0<��0��s�R�8��|3h�p*�]ދ�w�s�Ʈ2��F��ā���)Y@&�ON(������l��_��K� �Nu<k9��j��dQ��R ԧ/L�d?������5�����4ϞH�5����	E�y�AH�p����M7�����kd��m29?\L��y�*�`ұ����`�5�6?�:up�6R�1����T��2����#Ո ��3����;ݏa����3wV�w��d�	E�\�ib��#X����+�!��N�3ՙCZ�9-k�w��_n�s*cY�_�2Iy��{-��W�k��Nb�,�ӭ���(��%$1Il͘���yh� ��0%����|�tK�x���l�`rV!M� ���4��#�Ր�Wo`���(+�^�
��	/��ൾ?�\���bpYl�'B�b��g�O��ĵb��s2h��7l��/�S�R��o��}~��H���gG�v;2�j�4�zW��Y�f�DL,0�'I0�i��D�J)�0E�z�6��%�����7���~xi���!�>˛�S���ݶ��7�&���_d��|��O�L+o�~�����8�:I'҆�|�B��	7a���􏧜@0dx�v0��x8},i��=Z[�"(�{�� h�T�]�1-i�#�$�\��Hv�fR�������,bˆr�F��ƵCz�k�1�#�����C�:�}�M��릲��=��rx0���~��x>tR£!?����/l{ۨ/���n��T�69:f�|��H������U�j�ցU���'̌..����1��cVS��\b3Z6���n�\�f�پb���3\vC�N�{��� �ڨ%޳(�0j9�����h2�!����2�>|5Z׽�DFT[��8�~�X)@ą4������^�)6��]�J�^��=aH��í1��{0��ւs�;��-P5����9�.J��ȥt<����OKa���{>��L�����B#1񿆤�1'^�M{�TI��^@�ʤ���u�Og�d�L��6ht�_�Ý(�je�~������'���h�W����c��	p� ��
w����-�JL�����4c��lJ���z-���q�yP��>�f
(�(��sc� S�tr���2`T;�(Z�6����u�����ҤsS���tڪIì�Kb�x����)?v`��!c�!�z�sV��{�'g(��
Ll�N������;���㟕��϶=�"���1�e؄㄂�k}�ɦ�v�<#B�B�p��3�Y��~	F�{�!��\y��UR�脰]I�$7�y�U�]`[uz,����!|B~U�[Nn�f��Y�?č�}���W�頁�pї�%_�I�e�S�؃WC�A��LJ�R�!��\:�8&:�Rht�:<p4�Ñl�!w'~�A��A@3Ci���A���Y�d���RQ,���X`"�|�U^E�����K��Ō-��>��̉Ȓ7��/Cb*(MU4��4-+`��S�KB�x�=ûaT e�+m��$���0�ё�%A�6�m���P���5�M1���G&�!l��x�\t���pf
1����?V,�nKF#��ac��c���ԼF�<Zu���+P��`@�e�Z���,�Ȥ����C�cN��So��8�ļ
E'�h=��SW�W �ԕ�c_8�� X?HE�H�փ&����U��������� ��w|ڈs�ǧ��F���qK�|�Z��#g�/��uc{NL��ɔEmL�l߬?H'rav�$*U���tg`L�^�B�a,68�uh�*@TZ��l}#��'�8�j�4�Z8���[�Ro���'DM�̤�aQ�$��yL}��~��"��sx��2��ئ��DsX�GR�Z��p�<�r�5���l������Ǚ8����(����3Dឫ����f�F���������DN�Q_���!� <U;�����z#�e��N�n����.1��ܘx�@� �zm~l����u���Ҷ����C�������W�~w^_?�����)����?��������J��X`Wҩ��<��D�XR
� �$�?���5������>��P�4��Z�$+�s�'�C�~���ȋ�b��B�S)t ���'UJE��	�+,:A�3Α�ODy8O��o(��?7s8���\�u�Ps��jf�[�(�d+�]�̹s��^�E}p�����c߃+�
�
]18>��UV �n��)�J#���;ۈk�P��0Q�T��k>�e�\���ʭyzk�~y��f��2�NU�q��H۱?�ǻ�\�zFA� �#�Sh%R�^���ك(���'t3}����~�M�2�;�C��ЍZ`~���q
vy�ω�WR�T�6��<�9��p��������	�-�Hz ��{v��l�{���Nĵ�lߠy� n�|�3�k��H574'X(���/��/_�MU�Lo��Yt�cFB�~�R��U�\KӪ�Y'�h��odϣj?,���cPw�k<���آ�H�Y������'DI���'-}���b�1� �o�m� �5X�5q�����rp��e�F���o�'$e	!�֡&�F�x�`%��塀��<2`�V�F�+@�}l#:%&�h'�	�����H���"��M�^��B�x���I����:;^����.�6�o��&��ځ @�E�*F��L��4��|Y�	kz?�d0J������mO���\�w�#���!�b�{�bZ�<��6�m'>�;���|3����,����������^�M�-�rLTWV�@>���gq%6;���1�鷌G��~{��}{�r��/����_]i}O�������˪h��+�[�Ȟ��`QC�`d�|֢46���Y&{0�˦X����5�����O��E]����|��>t�]�؀Ѯ����N)�~m&�<����ƫ�Uu����F��㳰i\C�l2خ�9g�g&�yfC(G�ؖ2lw����܎*�s�ɹ��5�Cb���_g�fh���{ .*�3��A�@�q�/=����ec��,IP�¥����/9�����vt�8�ge�����H�h�нqZP��G��6<_E�b�ˋ�v�����al��X
(�X�<��Z�����ߓ)I^ɳsX�ߩU��q��}|͕��<��l�l�|R9�5P��z��@^�%�ɢ�l6�Dp���� �K��o�`6S����J�������������w+9_�i�:[��Mo&�84Lϔ��B ��莝��L0p�P��cq�����(����!j�K_2|�&�x�1ǀr�k�=B����ԉV��)�I���'�tn]F༣|�b"g�a�$pƢ��w�����bF��1�X�������3i�o�PF:�>˺D�y���ξnn|(�I�6]�������ob��S`1DMCwj�V�w{�������w��`��@�R39�u̢<�I�n���E@��r[�x���;��f{�u͋��'OF�D�xD|j��q���W����S��a����Q�!y���	-����-�A�<1��e`��{�k��f�=yk�Qg@�#�����t�Y�źm�.��Ӝ��Z;�cJQ�W��)k���n�?�s��������~��?���o����f�Y�E�߫��������=%�Ҕji���k[�	4<\����k2��PԮ�C.rhZ�LIw�.Vw���x��̓ӌ0�����w[���B@�I�t�@d㢀w!�
`�	����Cx�9�
���#>9�5�S�����K�Dst�z�j����$��՜���Q�#M��b��Z|X����ݡ���bi�
�Ւ��3v��'Ӱ��82)��O��7����X�O�T��=	�,|�ټ�R����uQ�Yz����+?��?����,ئ;��c������pEhq�$k&	������`F�����1ڶú���F��r�Gf����ֹ��/H��SG�ޙ�[��z��>t�y���o_-�뒱g�"bh�� ��<L^�u��x�Y�9��"�%����>mD�:M� �(���t�F�ԡ���VԥS�|XL1mԓ�
	FC�FD|fS���i��V�Sgq�I�k�BC)�����TJM�@E�M]��{�o�G�h�0I(EZ��i�|��!~C��:�f�[Cm=�au��yFW��'�i���>D�V�Im��������Ąe]^eq�6�������h!��ֺX�7&(��6�S�NV��#B�L�'f��QV�z)T��5�/j7V����Ku`�*�C��E�3C�Hyj
�8�3Dʦ��sJJ<7��uR��s�\Qn�ce���=q���=AJ�,�$�e�A
�A�d�����6;D����	a��?�H����t��咂�Zd��e|(o�����z���>�~�^n�Cc�Ϋ�d�t�c��ic��q�G'!���Df���nA{2��O�<�/�:�Qӟ�!����h�YR����PJ��\N�	�dn��ƔC�y��kEm���)�5�xI���?�R)V;Q�T�ƛ�MM���Ʋ��X5�'�t�Y�6D%��m/�ܫ;+0�s+k(M�ӝ!���QT"�Mg��gW��R:8��m��3N�/i6;|R����b� �Τ�Y%pX�3{ɞ+�tJ�'�7��~vW`�5+������wu�p�L-����)IH�{��3�+4�0�����@���#�[pZ��w����&TM�g
"��"��s���M��s��h�����q'�`@$��*ۓ����6Is��,??t=�kCZ<X|���,x �>S�z�κ.���	�I]��0`l��iH�yO��a�}�Ͽ�Q����3����U�5]��A��j$z����g�	�m}���X�`��YlՃ�m��zL�F�)h���6�z�\�:AH�6��6RxV����ߴ��$�`��� =l�8�{v#�G�f9�ًE��6���c�BQ�-x'SC¾=��esf��q����6����`a?&Q��] qx~�����^ʵ��m{Ĉs{��^��*�A��T6Rˀ���u�R�&�gp끵%����*k��ރ$�x��]�e�f5�aן��W�h�ݴ�d��:+����X�1�TV�QN9HA���G�xE09��+Q0X�AR���<`&���5E0 ������ټ	��	k� 8�?y��38���"`|����)ѼK�t_H��2��}��%G�N#c�R�����f'��yn�Oa���p|�����e��&���[w�d�/2�C}�T�ڭI�V����$��';�M>���斉1�V{M{�L�E{�iC�j�{6���������ٜ����fR�}
��f�^���5��#k\�BC�D"���E����,���߯��Qԙ������Rq)W�Sb<w����sHQ?(�<��F�S؇��C��\��mn9�����a���jT�I���,�>���S���O��1�msk]*��=�4s�yy��E��3p��R	�c��~E�&��i�<��(�����mq
�12�@2��m��a�1%��A0��r���=5�SC��f�>�U�~y"s6���b�D9�S�.F��Rn���O��2��{����婿<,�f��ﲒ�5��5��� K�r,6�|둦b�+���N#�#�M�#��f@-Dm�������`��?Q������̶u�O0���Y=����R�]�[�����s�#;S�͔���4���6[���F{�k��`�&� �a>�qm�KÙ���.f`b@��U��ã4=M7��M0N�*&�-��К�"�T��Q|��?�	#���c�-=۾�A���~�r��A�*�tnۜ5�8�?�N�Q>1����#(�";2�в+�?�dʕ���ӧ�E��(#�ˈ�� ��8�{�����b�[���m��������������w�<����bf�C�m�K��ŷ{+f="���2�!�S����)NWǱ��b+�}�t,�{35���F=��)�#��2[��VvВ�Ng�L�Թi��@J��W9�T<	�y�'e�":5U�']LK�r�:�g���_>�J�E�f2R�o�֎�@���x�d�g�~�2���|�03۞μ��v0�-�v!��^�!hH��� �г@�}�ڛ)��,�����m�_��#L�"�ߖ<~��b\I�Eu ����lǵ�o0�U�� ���cީ'cQ�5"��-<�k_�H�v|d�=ل�5��=T��s��^��p����6�����m��rdG��/�H�X�iB�B��͸欠���ˑj�VZ=�Hzx�h=��c��Y��4L�V��ؗɏ��g�����*���O���1�Rf�M�Ŕ�7�˂q������x r�m� ���gI6fMO`�kb���:�̴B���i�9Gl����9R��M��#�	�-5=�9�:'��?��ysie�O��A���qvh9����&�8y���)��Z����4�v���l܌ ��}|���2G���������O��-�y�zeP��]���a�9��5�8�m�>Ag>�?�C1�<k�,���IpQVr�%=�b�JȦ��D���2�cSw�v<�&陒�m��8�Cb����Lߊ.�6~Wg'�Q�Lh�J��8�n�o�6�P)yZ�)<D6��i/��c��!b�`A�4m}��ӿ�˿v���UK����}��b���O�ws����Q?S�W�!bI��CK:~��X��M��T��D!;� �~���4�__u�.zk�ɱ0��w@-�f���h��2��~]��r��T�S�����s&B������/(�T&�M�U�<��A;��Q2�r��Z�Bmf�6})���l����38��2�XA��e�e/��m��s�^�6&{��5g�~��V(��g��*����Vn�۫l���!2ӿ����0�U��z�v/vf��}a���O?������Ñt�}ͼ�ei��`����z�l�͸�r�b��o<��.����o�Y�o���3�c�|7.f��jiA�G��r�z���~��'��²�a,.�(�A���Q�2��Y��T����C�	�i�x ����y{�o���9��ß��u�d;D7�vsbi�O-�#�Qc����67�ӡ�L.s{�r�h���H'.1T��S�(Z������&�Jr����3�;
�	�F�.��g��=�4�f��ev:zШ|-L�>�
���u�\*��q�We^��4-��[��M�h�٤Ժ�<�4��=����'�9�'�P����n8+��KyzUY��d����6xt��བ)A�v��\r�~�%ؚc�dr����E����A�u�LCL�V4S��n��7� �� �f?4�Pf����8���{������`U�VsO1/3�D��J�,4��3�5��q~@EJ�X��`@���k������]��%*�
�������^X��p{� �.=�E���K�|�.]��J_|��̟��+N���ڀ���� ��ߦ�]\o���"1�'�?�\q�F�H!��)��y[�r���:�����7��f1K3�o�m��2,F�&6�15\���w�T4�cZ�ev�B�T���3�4#�4�2>���� g�l�1�����ހ�g��2A2-�2En�*�;��r�^&e����G��`W�%�"؂7�u|r%�l¿?�5���w�6f^�2�K��Rẗ́�p8g�d���_4?B�E��9|x�ٹa8�����>�ݙ�Ǟ�m�w��9�HA=�9P
������~���ФWB�
>�1-�V�1ŭ�s�]?��g�ُa�~){n��j�?hDb>E��ŀ�H���Q��.�+ ui�~��釿�!-�0!-�mӛ��ڔ͐�t
�e�l_�.�4Q�.e��'��$�	`G�����1�An��c1{���f��s��ߐ'�\�����D� D^k�n�)+c��9�f�0�8����|�_R%���;Z�M��S�.r�.����E@�0���и3uϧ��d�)ɘ��J��/�>���)l#�	 
#��v!4.�m��~��IL'�MV*�8�?�m8�����=���6�E�k���ӱ��2�#j�wŃ�`Xl5�$�������'>�ŭ[���Q�[Tr7k�l��\K��c@Y١�9/W�.��}qox�'����6��ujM�٫��8j��}/O�����a7��� ??�ǔq-�0���������������G�����G�Et^�
�F$ّ'������\#{S��C� C9�bщ-՜-���y;gm����QdYf4[�)A��G��Ƿ9�ϩ�8��̈Z���{ٺ��~�9g�_I"$Hp��y�N���"��U�u|��7Zl�AN.�)���a���q�Ћ ��,�}84En�3{:��њU`�{��B�8Z��r����QN�	�F()t6�'R�� /�2������V)71�!G�9踥��1�ߟ��zk3��q���/�W������s�(��{���T�"��_�*��7s;,4�pMYkw�	�͒�%�g5a+E���e�*+�_~���zh(���1�z���q�(���J��-Y ����Ã�Z��b���j!D��أ�uS
/�ӧ���]ş��t���iX��e��.W��P�2|��N����:�Z�}?�Fܰ�H)"j��wD`Ҟ�h�X�Ŭ���1:1<�z���o�����ĳi9[d�Z��|o���1)�N�B�m!�G%��8-���0N���^~	\'E�)��?����i&����[
�1�kV���GJ�Y�,����y}���:L~�݊�?��O'K��H�#���l�>_��5#~�E2~��c�C��&��@C"����kݚ"� ����xP�q]_�����!7e̠�����f��iZM�
d��R� �' ����l�$V��<e��0]Zqe��c	մ�*�cyN9 ��(<C%�������lB�]�6����=����_�o�_DFJi�����lS��oI���I<����`�9��$y����Js�()�(�����@2��� e]�H.q���@��� 5Nf�M�`�#�X�$�D��OL�R�
(�Ȟ�Ƹ�h�XY������~8)�A�q�OA,����6���ћ?r�&o�l��9b�X�\J���kQ{56���Dyb"�;!��3��o�G����=ci�%��B�)�J��YB����%ih.��io��amE��EU�l�3��٩��(��j�p uF�Ns�fLў=�{��i��?gh ��{��gs\���C����p��u����3�!r`"W���.�'���q��٭Iz�Ơ���@�����6�|���l9�	Y}I� �����p�gl��#�+�m�/_�87*N<Y[I>���OZ��Y	�����˛��uL�Zln�\��0�-Y���PO�o�9
��,Q��F��w���(���*SSV=e�u�<"��fD����ʹ,�]o�I�$���Gd&��ۙ]�-���H�����_��[��},yw�Ù�* ���0U5� �����F����fj�j���q��`3r�t�\p]i����3\��AȎ���˸��CA-�M��yژ�*2 ��@���
��zG h�� qp���SB��MX���=�I��2˅��ޡ}6:X]�nҁp��:C ���@��z�d��hR��~R��4��h�CF�ó�U�F=mN.��d���L�'xI\���
�sq]������w`Ls�ac�[A�qL`���B?�LPm�^?�U���N�CI*2
�JURt�ܘ>�p�*�
����9i*L�(f�0/RV�����R0��~dRa읞��oǂx��Qb����>��ׯ��~s܄����8I*ޘB!�-����0-	ucQ&@)	1F�dJlL�R���ͳѦM�@�"&ؑ��3�}z�j�5�spnA2a&BH�_H��u&�p �o�f�2�%:�L�Z�$���#�%uZj�6]�Hq5�;Ʀ��8��pwf�}�hB������V w(,��Y2
�z�i97�8�L��.\%�{?q��z�g�*[��	��mH�{2�I���bB��h���	��Z�k�#��˔��� ��%�X�Ue_�G{'�4���[��뮟a�O�F�|�z�!.ɂ�2�2���mEݎ̮&=�%*�/.�l3:����6<NHt��p]���;�'�G�WCe&GV뮍���_�aI�(����W_7:hQdT�jt-d��%�R�����ww�����.'y�O���M��k�׷7�]�����~�7|��c�"�Z�86�(�b��ȹ��ȣY%�Q�S5u)�Nl;�8���+��:y��_�,G��x�fΟ���DǙԑ�{ʖt��/1�~f�f˲0��.�9#�Oók@��:i\O�w6��J{d	݊0�9:8o�t�����պ++,�L���;>���'�Q�<�qc7�`��ĕ��ƃC�|`��"�GFQ_�8�����L��І4��{V=͸r�C������D<WB�_�+��@\Od)�^���/�^���Ab+8����"]��v|����l��(�,�33�����ef��|�3�w��Wr|�>���T�|js6Z�+�"XV���Ɣ3���~��p�///v]/GD�FN�n�#�$��]���gE�F:/���Í���	G-R�����b$� �b�\��%^_�Q��U`kW
d�5�k셷H�#�=��M����S�?���'	J��:k���=Iu|Wc��UK�A��h`#��@�m�L�ck��; ��G�u'R���%�_�=Μl��Z��[������rl\��^i��t���=�{�]��g�$����s3��cv���,3��4.%4#fA͆v��YJ���xN�N��I;�G*?JQ�1=;SfNe�w�s ~hr��U=��l�x���(w�U��]l8�Ճ5�%���?�F�E� �4�|;v����	 Ab�_rB|�D Ϭ��Vg�Q���p�bwfrl/�Dwc6��%�� �=m4���ƅN��̮�j���\)#��|��4e6�k�&����M�'_N�)�U��I���j�D���i@��0`)VOAtn�dC
��9;�vey�,��MA�\��"����YL ����M;��$��	va��TV��_W�M�	?ݛ(�t"�����,M%c^���6�`
݅u䑩�b9T�O@�zH$f_)�x���^���*ƭ�|f�}^ϻ���2롳����7�я��1�AY�|���n>͘>��LIy��7�e=�{cFU����_�^m�01C2 ��#?
�(?�|�ƃ���T���b�FK�B,�c^r�*�If��>�t�F8�u=!Á���Okf������7��o��o~;�n�hH���8������k�|�I?(������6n�����z}�����p7')�����̖��(nj�pOp3+��*����Oڗ7.�."�`\��P��S Ԕ*]/�r�$>gUf���H8���ASɒ�`#H����*~_�Ch/��ZO4�9V1(�ID)~��5]"^�C�X.�V�ˤ<�l\�c�j����� a&oG� ���XIN���IQv���0��]�V��GO�3���5>�.<�-�utx���l���Yצ��W֠"�͛LR�l��/��a�p��"�۞)�����ʜ2��A`��36ឞx�M�����0��C��G$�2��i�_5
<��=����DQ(y�;��_� �\`ｷ�ս�@U[R��$�B$�J�8D�����HD�)S�\|F3�oJux 
@��a��-��FJ��s��I�,�(ͣ�*G���F��.4D�Ԯ�$�@����k-r~�e�֜����aG�HԈ)��6 ^�����F�ϙ��_��lb��'LW �x��~��f�Om�K�b'�Ic�Ñk��'ep�6��Vb�c1�](���3	+ys8e��.�L���g�g��!�f�Ό���ڐ��Y��2�k_,�(O٩W@M�duxg��hR.��<T���R�Ф��3�<ܿ� �g$D�|,Ȱ���m��PD{@)��P�d	?St��B�%�W�"$�u�Sq�xÓ�N?�ݨ�`��:�
��h��9 xm���$^���(��r�+�Ck��F5M+�7�T~�  �IDATj��O����Z��>>v1	��颋�`8ҳ6���L�@h�æǦ��-	p˱a��Q+�Ү[�!P�%��0& 'i&�ܷM��zƨ�1T7�����+%I�,U�?�b�m$4�t�7Y���1�CI�9x����@�|���G�F=[:N��t/&>8#��z�2h`�����7���,���YXR
�Y*����Z�l�j����l�{��2>F޷aj�ڻO�'��#�n��$���,�5~�O����`a�LNہ�`�H!
�p��t9���.��e���9�D-��C˘�ǘˍ{�C��q� �e���厖�^w��i�AW�0���N������O��)Lқ�~)$�5�"�|����hq":�U�?������AAkV���>c݃WJ$~	=��\�\�s�ӳiB8W+�DF�cP�#����r�uަ�� ݏ9ScVVk)�A�@Igؔ�AN�-l%h����d|����ޫ�Oڳ�n�D

K99~;�<@�d�!�T2�tRF�V�:h������6���Ts�\�}J�:e�3gͱа��'Ld�c mX́��B������S�qm|$�{�"�Jl����]�1��~�[tJ����k-e]_ �82F	89֮ =�f���Z�lɃ��O���#�f��l,p/iLd����8������{@���,�b�i�����x�z���eF����2&����7�$Y.���ܻ�z��isWte�􌔈I�=�  ��bܘ��pC`�����@X��ŠPH]��t�������M58-�Rg�ٵ�/��T�� 0	�R��k���ղʀ&u�: ?Q��������"���PLvf��u?Z���#N��ٕ�ս3�_��CY��0ǒ`��>7�_Î���K�O-y�5�R��<G݁����ѭ"(Ma]��\�j��;��3-����L�	@��%G��U���Ƴ�&��� E�|_���������#�A�As���ԯ�s~��:�Z)2�!�zo�h"�zjk�Y�A�� F9������q�R_P��h�Kk}����w�����M:���Zi ������J��D�,X�&�K���d��%��v�m(���*pGP�Ww-�~d����}����G���Uˑ{�`Ѥ's�e��8���3nl��h���'��M0H	��c�m
7f%s1�2h}X��$� �%�7�ڙ�V�x�x�2�����W��H;��HG��[�z���{�ܙ�O�}fW�}Tte�Qx��� L��3��DM��%y�^�$۴��(�g��D�b�r����u��M���m�I��a��ݻ��>�F)�� �L�}��9vA惡l�e��ȘR�@���6 S�c��2%� t����$�[�/.L�kn޻*��29��l�(��u�}�����w�*n��k����c ��Q��EP�� �5}Ey��Rܑ�Ƥ2�?<[=�$�Sɪ��,��e����;�B�4)L�r�'�9Q�9��8~��g�����ĕ�������nRNqz�DT�n�3���+{�1��@hb���t��;TfҋQ9Q��UFDg%l�0���Hk1�rMM�6f/��S�A�q��|Y�N�Sv7�&��,"�cs�G�4����3� ̘w�8x�Q{O��S6���4%�f�����H��[�����46Z\'t2�o��� ��.�MYSF	����f��}��{]%1$O�S�����,�(�yb��KA�$��$aK'K���΢�b	�Ӿ�}�<�d
#�D�] J��n:�h�(T
����"'�L�/�ݑ%�����3��A,�p
5�z�AΕ���`�}��ܘ��X�2�9��J�[qI�|��d?��g��D]�^�%�"B�l�u��_�uv�"<q�r��P�'M�� Y�����b��bZ�Dsy���1c鑍t�[�Ɲ��o�/ZO=[��,���uuS6�#�����~̌%O�sh�aS�h��$��8�m�=jͥm�� �^)X5�K��(o¯ ������b	Q�ܐ�5��u���oBO��\�y����4rxjAJit.�<����vx���q�@n��AM�-Kr0lܷi����'�g��o�}��������6���3��A��{�'JA �C�;�l_��ZC��NƼt��Zgg�+��c��ڵY{��`d��2����i�##��QA�|���3�K�,��X�켴��?I��8\6z �|���=��[����/��G�f��C}��I�|�^��
�2&3�M�f�c���x�ԃNSf�-�Ok�7g�F6�@���:�#�/���Jp)-nv�����S������������uks1<���������*(L�����mpl4�/+S����4kw����Oy�L�$�a��Ȉ����7��'ۇ���L�ٝ�SU�H �2G�L������]���i����αQ$��/���2��G��N�k��)��i +��R~��l�˟�����D� <���k�tI�/W;v�F��h��V4�b���:2P�zb�Ɛ��H�='����3��cL�wA� Wy��khR�Y;?��Hn�yI�۰�KA>��'�=y�>�sz�Ï?������}Y��!SS���G7B��g��hw�</���I�.t��|p0�A�ל^��m�S#���� <������1����E^�[ᙀ���3&�:?�"sc���;��:�m0�\�a���0��"1�_�NG;א;js�x�PO6�Y�.C���/N�}�l��#�LxO':�c'�����|�kP�6jo��5ةQY�R�s�#4 E�b!�z<���&�3�t@�f�i+��1��Iٯ� �_�p��:]�	n
1`�ԙ�>��n�z�2v�$�Ko�D�����^6"�.��K�B72�6�a�RS+?�w��o��\�l0��ܠ\�D#�U�ue� !��/����x����D�eɖ����Z8\���>���.����^(P�B�ձ�2(��:��<��+�+c�s�0鷏T��ă��e�:�Αd���p�RPy��3�3:�V�ehC�yU���=���܏��E��c�\�Y�؞��C� �	P�aw�)�E�����&�b�&����c� ��� {��=��-H?�;�`���&~EK"���QHԢtY�L.D~��Wg����U�,Otg��q�l����">M����|%��,[���a��f`*/�]H�j���m�)��ޤ������DI)�	`(�
�yZ�ߐ�7�2��G�B�+�U�0r���2G�D��=�R2���/�)�Ԧ�(�D���nϤ^�� G�^3v����3X�5���m�Ojc������.��i���6z ��T�+����J?��,o���$��{���?ۿ����+���������fS ����� JR�Q�6�f
L��Q�χz�M8fo�Mm��)gGj���z ��P�����=�%��=�EQ����6�#�I�5�b��@����c���~i�fK
�s���x� �Ebsy��,1��F-���+�v�%���� ���:��6f2%|?���p�r����n�G�K:�F'��à
�=cg�o�z�艁����XО�r��/5�D���n�!���U���э���У��m#I)2���
Z�&�X�"n��)*�#�B��/w��k�=�,��`���oN������>��w�MTG�4:c���N�YD�t.n����+]"pOj��&�\F7��p7�傾�ž}��0�^n<9����i��X�� �6�96�M�k+7��e1�S(L��)W0��3m�J��P�5�J@��Y�i'jSeT����e�K�wE�- AF�bT�z.���Vz����i 8�nb��%�Q���c�R+��t>��k�B/�.q�~TZ�(\�_����� ���������gFwLO'��v��l�ag2�݈�]����R�bJI�n�8��_���� BD-:U�p��~F	��
?��6nrEl����Tp+;P���V�E��>F'�;�P�����b<K�<���a��D)��S����Y���ԥJ��G���p��O'o�uP��"1C�?�1̩���2��� sZ�o�wlNҢ����:�Δe���cV���u�E��3O8
�.���*սY���7�O�~����X�aPRl��M56#�ԏ��&����ɹ��V��Дi���o�E�Cނ#X����ԍ���M_/���Im����%�ݩ����[� )ldC�;^��'A6K�)�M�EQ�9Og'v�"ۂ��Z����?��N~��%��X��c�)��!��P{�|Pv`�����Q�G��L)~"`�bJ���\\�e��{Y���s��.�M,x9���\ĕ���{\//����ΦҊk.fH�����{|G��#�L��Q���_��.�����~EI�չ�VwS��g?(����#�����'Y0�U�4d	���l��z4� �����$�W��8T!F�=��,�N�q�Ggxd�ne�ٔ?�g,~�\����F���Cm�_;U277��@"� �&�^�'�������@���]�wԏ!>!��_��&md�@>�]���0	;[�Q�G�:��]���,څ��-W<��JA�!/�
��{ ����Ma��w4d��5�>|
FnxI���9	V�^6���>R_����!8bނ��y,r~b�g�L��g��.�j,�Qc������y���5E�ݑ
�r�kߪI0�J�,�mT��/��.��׾0��s+Ȁ:ft܈6�s;�s���\�䀴m6�q]��+�eX�kV�H0�A�?�*�<0�qM!!7nrh�$��6���w���!1�U��Yo��;�&Ht�L ��8���븷���������O��A1UY��Su{P��Ĥ���d��@�hU|#x,?�Y~Ҏ�a�>j9�>�Al�M	E_`@��F�
x�Y�PZ�6ش��Ë4+���I 
9t.�x� �B���v��<!S�7E��\��6� ���b�D����^|�X�@ﲼ���)�aG^����/8�$������-ц��Q���#�@����B��	�û���F5�Fp8�T������I����Q������'z	��N2]��n��~��S-�ǆR�������%[<z��D�n�p����Z�~��|���Oy/h�潌���zl<������I}X�NǴ5&����^�^S�y�p7��l�n���,��b*x|��>��p��U~��؏�������^�q�l�,�]Ҧ�8A�^�G���a�����*�$��a^,�SH_��|�3����=St=l��9� y��d�g��6۰��=�t*"�Ī�*��0"m��4n7�SX ���7�b�p�X��AF��$?����
�Mz�=! 0h����LJ6}&��h�v���y.�۟��>�sE�UD���Uedo!$�<,2ݗ��K4r���q���&����Gi���S	jbL��+@0	a�א��)��?^��O��6X�暚Д�xM��<��q̟��L��	�rH�^a�ҳ�/�
�X�k>lL��<ù놙)�$�+����u}Yn�r}��ҡ���A?�L�^��~������X�,�j�@����{>?_����X��u=����^߿�S}�)E{�8�m���ѯ�͐烑���`1��G=�Hv����T�^J��p':!�zI���?�n_8�7�d�&���5b��A���Y5	t�)b��[��\Y�9��פ~�c����<J�n���P)�����u����������y#ۼ��w���^L���]��*���ʎ/�0q��	�NZ��Ub�EJ>3���9Oәq�]��C�e���u���T]G���sޤ�w[/����a7+�E39Z��U���s{&��P�ե`�}�6i���ܡ��O��Yd>�a?hӸ�C晉cS 3˶ą�C�3�*7(���"��э�8�P�<`��������ք	��NA\l�tz���FR+U��ž~������)�[ Lx�ιE��JN \��L]~�+��nw�l]��!��4�ă�����Q[�6\=�7�a7-���F{�ky��IG�Yw�qh�_ΡY�"Om!�}����M3)�fc���m�7LF0:]N?�w5E!2`i_��׫E�s��(����ܐ�ߺ8ԾA��.GLrO�����Ó�Q�T����D���me~�� 1?f��w��/fF�t7Vҋ��Ӈt�L�=uI�&�aѮM\?�kq��2�ӱ/P�r6��(����l����Q��S�?w9q��Gw��@��I�ӤÃ�O-n8�+�K����E���d�/��r�JF�7�֏�$ ��@5g���^z�_n������~�Jk�? e�5�hA��қ$�=%�*�R�B�����@̰���qP�2}5e��9M�1Z�H���䪖ӈ���w^bY-I�?�G b�Y���'=PJlI���zV��jA	��e
o�A�Tnvnސ^���_�1���3�5i��-�u�Ȱ�dCw�<R*�gReGO�
�Ӵc�p$�����3ǭ�����"Jqu����Iq��DweF�),9%E-P:$�4�LS�g��ejV��2|R�2���=��oVa�V5�O�o�:pY�s�m}+��m�O#`>M~Û��W��h0DZ4�\������#;0�Of�D�I&m��c�b.ڄ��m�e��y�(o�г|�>7��C��Y�ӭ�gb�u7>�����b?��3N*���ʴy�8�Qoٻh���������hy��s!	h�c���Oق�����`�C�����H�*j�7�IehEF����-��!9Xv��T��ب�/@f�L�����;�0�y��������� �����qzzWj/����Ch:��F�#�E:�nk�&F!���7�Qx��Mē�ӥ��ԍ�O9�m�p���,OXO��](t���C����u�������'�����U�����+�7_5�oq~Md	�Zu�r�ۗ'>3&�Ыt�f� �e�O ���0s{E��<�������)�J�"��	��T�tI��w��M�����)��`�M"=��Q�u|�3�w��=y����+ ����#'�e��zc���(���^�%���������l������h5�|z�B������=վ���O�^v��WX0y׳}���w�CL���7�Q�� 1���
1�c	�����A�Fm~����-jf�0v.�(;�%N`β��E�Ȟ���h���:�R�>l��
kc���m�+� ��0
����9���цf%�ə�QR��b/���:]��Ϲ������?������x�L�q[����8�"&q��&���񺧘h�i�p�q�ojY2[r�YQq"�/�Y�
_˫���@��cU�d���[@w�7Mq��*���E �Ć������M�Xb-P/vM^O�Up���P�T6�υ���Ȓ6:n9} ��v9z:�l|Vn��;��lVl�d�!���DiKnDt�x�e�#Ako|�&w/�W̸1��ڷ���z_�|`�Xxމ�����~�W#��{0�{��D6b���i�zl��E���}
(��?�d���� "	#P��%�}i��t��R;��=Ԧ�O��g��)6H���x�H��2@F  ՜�ȃ�|��5��<�{����u���B��/ �3(���dp�J:��ض�6K�=�>���庉e�һ�����p�5&�l 8������	w�1�L0�Op�w���.|�4\���=kX2�vL*��}6��`�J���#J��Țx��Bt���?=(ݷ�"pV�0$A�ڐ)�D���9�p� 1D�!s���T�&2�����˕)�o��ym5��S���+�I]��]���*p�r��ͼ/ ����p���b��<?�d������?�����p�I�>jE��΋�#�5�7GW��)9���O>�P��EZ��2|d�)�zn���k��X�����9�Z2V��aG7���?Ou2"����"��T&�uFy�Y�8��eQ�d�>���^�h�2p�=�|Ai��+X�I]��!�f'%�4VA&��ɽ�8�T�����3p6���MA���ka	D�WQ�ġXc$C�	<[�  B����̫԰���#Yό��Ƚ+���ۮ��� p��vT�.�en�S{�Y�$����5�ċ��@:; ���y�6�Sٲ;D��K֯���N�"vl%BI?Y���+���:��'~H�g,)<9�ǲ�")O��0/>~�Ӻq_׋?\oy������������ ��YNdb�� gl��/���>n�@��w�$)�����`�d=J�Y"��G���&�"�����>H:��Y�t��`&j�&�<�6�ae<�������,Lt�^8o����F0V�� �:����g�1�;Km_�/��uq0���<�b��I'jẗd��1���W������_�w�[�� �g@u���/�/x�\;J���`�� ϩݝ�wfH�f> [�����u��-3+�7��{�d�tܢ�dc�&�(�=J
n�,#��ΛyHGȨUft�0�Ckk��������r�����$p�@W�	��d����hx�����3���V��P�Jo���v<�U�>�G)��?H`D���y�i�+ҟ�9�PN��=^^^�?�����=�8,�LҜ��ň����%��k_qrc�7��q�±��G�qa���DV�V��k�*n^o`(��nP�6�m�<7�2�	' �UmI�����&��	1�Ɛ�,�"@ 1ˆ� ��Q,�NH�,\Q8��W�)�7G#��q"�������R�󐃺�ܜ0�����q�o�ڝ�Y�zw�N� j��mt�EsW#�iT/�e٘���ha��@��7<=c�H	�Bj>�����x2���l�r=���F�K�ZS�S�-Z3V;2t2Nc��0ܝ��P+�8=)���U��<��+yf�~B��.9�J��q�H�����<��,0E�B��gu�܇���H����q��������~���QTl�����ZM�S�nL��GlLW�xx��K�^wW�=�t�ٝP�.H�9gb�C��J5/Q�s���b�.Ys�i�Z�x�E�.�!��l`�@��xm�]�O i5e>�| �9c�������Y<�Q�4���G	wn_`%�U�E���6u�A[�3J.t�,�}�䥠-f�Ր�у�/�K���ݦ�:�(���?���iW��bE ��L[7�t��)�R|^S
ٿ�6B@����r���S�]��5]�0���C�`����-
,W���F;O��av�f�+z�I���`(��{w���U���y{A�����"��X�+��dQqg�V��'˄�F?�1G��~Hb�	;;I�T6�i�#����2�	\ݍ9�4d�Z�� R� Q�w��>s�������������¹\�܄�
4�p��L�؀�cq�%X�~1g(��\�F���ݶw:톾a��;O��	�I&i)[x9T�U9@�P0�)�����I��L����-;q�i.JB#/2�m;�{'S�54�}������2@Uʚ�t��,5��#c��t�>:�o�DqS&W���4A�����(�ڜ.��ھ��h' ��W=��k�� ��Es��nʄ�#�-Y&����Y)�t_5'E'�>��_`�M�q���g�Wn�tA�0�;�����Yp��$zGP�����o�`���훇T�0v���i"1�F��Q�A�K4��2� ��Ӕ0���tc��`%���('O�E$-�,�0�Q}��s�,�(N�P���.���?�d��o~PV� ;���}�&���N�_����en򮬂�,$���5��B9�@O6z�i�9'� �$�ō����R@]��F������������v�6���jeƀv]ʃ�U[��HV{�	��'��X�fa�d?�Q��y����R�P��i=S�������ңU��������B��R~k}âX)�[���3$��_̽�
:̰���8v��%���`5^ԭ��H�}R��C����gSv:qF�L�D+(7�C��V��Op���q��6��{�������)�۔)x�{�|1��D��~���@Ǧ���pЀ�f��4l��o��v��hx��m�Ƶ�E�W�Y��&��0
�����	�pO�}e���|�XM�8Z�Zd��w(,�F�de�d�v��>�d�b���~���2��l_~�
���e��@�g���&�"�/遲��4�xb���4����E�/��&��ȱgޗ�,�SN��zף�t�.q��.ur�X�F-k<�Yo�~5#F�Ƀ!+���ˀ�'Oӹ��h�&Φ�%�E�nH��qe������L�	`n��+���g��[�͛�p0�Vu^�p��*�0��:���Rɳ!�H������,!���2q��z���In�*gu��ΈKr�"�u>%joY�u���la�H1�fׄ8���դ���!��m>�]z�B�	���05GHl%��lF3�y|r�29�/��q���,��j1q<Y�ǜG5 �	h�3C��3�"K,�o߾�o��ٔ"�~�_���V-Z����ѓ5Fr�s�*���4S*@��E��^ ����՚�&)3�\K���#����,H���{������B�aE�FR���m����'��-F��z}���"��2;�gdDcx/��L�.Q��5ۉR��q�������ѫ�щ�}�'ވ/��6X���6g�e��`�~��tM�p����!�y��m���� �Y���v�N��ό@�0��d]0]LR~z+��d��Y�yV\0\zG	�!K�ً��_���h%9, �Ng#���Ji ��)x��15�U��&
ѹJ���VU��a����_eg��C'x쀈�r쓒��eV��� >8uM��6��Y䜰C�"��g�;��7��U�pϷ/�Lf���k�w�}���ۏ>��������/*m���׆��HL�b��6�d�3kQh��zEE��k��\��iǍ`+��Ӯ'p��iY��{JP��1Ж�i�����gm���3H�����T�}l��򹱜�J⮖xha#��RS0GT:��H*�Jq�u9�ٜ�Ğ=��$�Vf,Ne�G��]a!2�^("Z�m���+0u:%ѻ]U��p��^������\k�M��I8�E��q��u~5��f��3�˱����w���=.�2!��*�����v�rLܾ6������{��
N[ӱ8��;Nr<�-8#=���Q_��x�s��c����ǽ�=$�2���et+�*4G�zAGm]��ո� �{]��<��A9�1~9⯚�|�2�����L���=]	@�>P_�8�>�F�#�ܟ�\g	`�,����G8�`��p��"sqĄc���o�z�uw�n�\�O���HJi�� �^���s��^O�wQ�q-8ق��d�!�Ei��ф	0���*�3!��`�z�?���(f�9}d�/T[�c�P��Qޙ�rʢ$H��݄��Gh�B�d�]��(u��Ƽ��Ó�������u5�R�]<�S�ttI����u�_~�������zZ��s�B�-��p�V��\��<?3ی���]|��ڥD�N��w��D���)Ml�)�� F�o��BkCd�p�׀�-Z˨MĢm(� �����u�&�C.��K�!�s�:�=��$�����#~��]	�����zՃD��i}�n>�V�\Y��L7�k]�B"�d�V&@&(�)�GΩØ���Id'tC��C��L���p�#t}�𦀯_�澞��t�.�oGg��<�f�.U��q���:�.`L�_��	���c��FmM�`����&��9X7S��Zs���k����_�#�����}ٔ�Tl0��D��k�W �K��gY�k�}�3m��i��q��z��df9!�2c�1ɭ���LɫR{�\���la���L���<���0�?�{֓ }`U�d&;}ӚHpעz��'QNm�N"�o������@�"U&d�6�9:�����(A߹*׼�CoR�-/��c^p��C�S�X�n��s�M�?�zq�iH//�����ۥ�E.P�בV��梧�$�99���A���؝�Ȝ��.�ߎ6ic
�^U�H:��c��Z��O�I�MtV��P���������HE�^ U�~�#L��a!��#�3x�-6��a�bb&f�}�rA���V�c�"ʴ�_�8aT����<��|ȻY��%0��/F��e�������xjc~0v �v�g̻��m��A���}T�F� ٩�m�"��H����o�5bpm�����xQ7�}'���QP��r�0��}�W�~�u�.Q�1�L�q�9��g�e�{�����) `���2�(�`�JJ�'�.�������tȴ�E�|��-�,ǻ��r���l�wODT끃4���;���� Je��5�������?����/��Ͽ�r[I��)Z���3j���GD�H��X6�f� V&Wn�鑈��]�O=<�B�'H"S3�5<�,ov�YJ�+u�Oj���A:R<ozErGj=�t�`J�Af��?�EOeV �$�#�s����dYLPe�|&�w�G�?J�de5��ݯ�3]F�Ƞ=;�X�2 6rpJ�>-6:7��$m���xm`4�O覱�P�+z��5���{?�R��3��9���0�`�b�j6	��Ņ̮��h�`�z����3���{*�B�����.�9��gV\"�X���2��Y�V�!`�/Q��Uo���V{Q	8��|B��3��S�Xpx�wJ���9��܇�=A�K����+����Z�el����Y<6�Q�ro&^������O�7���o~��P�w
@K:?4�N͠��&Xeڌ[�X��T����<�o�;Op��^�9����`PKhZ���m,f�$�[��3�0�uN��=���{�&�=���"�kGX��C6���vJ���Um�������/��p�/��pSs�-՞�z����i.�\�U��YYD"Y�E��L�ӽ�N�B���9��Qs�{�����,)&��Pg��ߌX�Uje�^.�):�^�"�`[Q���y�S��յ���������L��E���Yc�J5��u���U1C59-�4D	�a�x!&P�c�ű��+��&ߎ��3:�	Z��N�������˗��`��w��_��Ҋ�Iق���������}]�ٽ3qx
���5�8�Z.��P���� Q�&jv����m��Z-,�o�he��3i-��#ay}}����� x�=���DZ�o�c#� ���]m.
X�>\N�`�@R� ���S�9��Tq ��b��Q�*�M�e��9%�qE>����m�KB��z���D��hF��}���v�N�:��7��4��R�`�3��Ȝ%����p�@�ЂX'�N�[}�X<7`$�|T���['�rR����h� �Y'.�!<I�7]�����"}P�bD���P��7�_�'�8�]!�g_~����a�QZ��k�p4�3u#-�<��V�����@�P����al��$�|�a�S7���?x���/ s�9n��"�uj\6P 8���L}F������P)s��}�k�b��a����h���i���V+���4%ߧ.��bR�bĢd�tC��@8�Ѕ�.�i����z��?����^�w2����)�?��T�Y'E�_�*��Ք���4]����M�`�y�dlC5��L��M7����Qk���.��+�~���p�뽒��]ˠ4�EF�x �͇�/��N�`'R������k�9���������/�+�Ȑ����6x�q�gav�V�B��$��Y!U�l5�V�e�$`͓��@��������"��/��T�7��Z�t�<���A-��:�KJu1�`n�,�L�IE�k���{�:DT�Npt�6l�����(���x�!Ly��a5H�T�cȒDP�q����\e)��0��I5t��KK���Z��hd�==��9�i�����^,��b2������O'�0�fee�U
�켓B��ɒ:
�=s�ӭ��u���}�|�`�e��~�����m�LE�]�������<n��9�0Nd�.g���G>��ުq�C��������s%�m��(1;��`w|N���Q����z-�dTR��G��[x26���ѳ�L�`��-Z���p�w�S��&mHI}瑻��/@#ȋ�܂�Z���v�h�Y|r�S�Ü�^�1'"�fS��������'�%d�G�u�U�S'"Ր@�\$+�P�q����Ȗ�dz֜\�â��
1<Yn�m�')q-p|~id�dE��ZHu��`�<O�}�� ��1���IwZ��Gx������%����Df��փm�6��5��"��I�N��]��p�v������ޜp4�nR��Ұ�:�P��@�D0ǆ�E��,otY���W�q��ˑ,x���o�������_]�ԚssR�8��18�8�W?=k%�7e<�$σϻ�W=���� Ȓ`nP�a3Ef�����Cd2��g��=N���������BC�͔-<�3 E6�|~��o��}|4zk������%l^�b�5i�@Ѡ���g%l�F]������tu�\NA���4\��~�}s��-�o�X;O��?�]��i�A@s��[�1���Ѓ��,l�K����0y�M�;׋�30��3B٧��Y�e�H��g��3�d&�׾ˣ��y�R01���L�����s�{��`֢2PeY���Uf)}����"÷ѯ�O���t�`46鉒Y�"xyAT�@��`}=�3}ԗ8t��,v?J��3��#:�ѵJ���Y��d >Nt�t�{������~����Ηb?]~s,�M��"����%�L�	��H��i�)�J13O[�'�rw��L�����Ӌ9 K��x_�p3�}�.À36�f;��^�<�����R�7�h�ah�a��Q[��ȃm>}PFdg�qNd�� R�)�`�p|� �`��e����P��ILU_,�-2��D�b��?(<bK��%�bF]J�Ȇ��3��6��̨Ԋ�tw�P��ɣ1Z~IA�	ό��\:$9��p"�ETJ�ǉ\�@m�J�
�������uu���=��+`'pl��,��2Ղ��'��d>[e��#��T�����e��X+�����k#�L :��E:l�bU�AN�x+,�:��P��m�s���S��#A��\��Y��33J�^�<P�fa���޸o�3�{���;���IO����_��~����sx�: �̉�eD�r��-5ԶY
K��2X��K��d�n��
�Ytjr�;�9)��e�r��&��;@WRԎ��,!�hk����sJug��s8�h��tW}��RHx�a�����[y,�Ü$1]�cp��H�+��&�� {�J�\'gi��cQ�:vf_�(�s����2j��t�Ƅ�\w�L]_`:E��% �������
`����+�ΓE���gha
Cs\N�j#;
̆���5�V�_�Ϙ0T�Jئ��t9���	K!l]���� @�!+�4y�'��������@����b�:g���ۇ��_������ �Pq����Ueq�U�f�?c*�P[p}�U^Dƒ(t��b�F� ���|d.��nS�x;��qz��]����@��m����k�d&v9�iU#m��j�f�Ú�w"ޑ��7� Ȣ$wYhu�\ȕ�f���rBUsCS�i�'J�渲6����m�DAW�[Z��ۘ�	������>6������y�Yw�S�3�G͖��_����D.��s���:��a�d��i	<����؉;�������۾9��X�9��+O���
�����x�>^3ڼ�E`��F�8��_;�P�y��d<u��]#qB�������v�d �:YC���-	P�3�N�RY&���1uЎ��xDC�x���VG��t�I~Ɩ����=�ȭ������Oa��+)���ɜ�ʓ�"t��na����82��A�����a0s#���˟_�������7��������~�W?�/�A.A ��A&y�����na)ۮD *H�买�������U|t��A?1e2S� kr{.>�%m�97oBM&!�^Gpي�������ʍ�H�ô��7���IC~
\]J��&�/�������t�1���ɞ4jdB�!?DI��9˵�fD�I�V)(����=����"��ώ48)��B���0�M'����z8��T)a����;ǽy}������jo�wJ�;u,��>'}#�Q�_���_�-h��VA�B~�1��|%8�@�˅�n4���G�Z�T���.�?|�%��y~���Ӕ�����KHgm:!�c\����ɫJB�0�� ��a�ߕG����Qμ�?�C���l�*�7sV�w ����,����;p���>��mm�8�	rF���O���No�81���o����_��1<��_���7.]��O���I�!�4'!�i���LO<:7F߂��7�E�crL�~v�a��8�rI�DѥO�3ޝ���jϢO\�Qe'��C=d�E4T1GQ8I�6�z@�8��B4�I3�R��1y����4���G6?�wF���!W�ǘ� �3��Y��Hޖ�X�,ٕj��Kj�͓�ܵ���}��q,H�(��pd xV�^�y=��pȖ�6�;�,�߿��ɒ-��x�p܎���g=��iw�3��fdЙ:��Н�I"�rN��<pY���$�,{��k�h��U����rv��u�'�Y�Z�)�O��?[�A���nd@y΍��˪}ٽ\ՂN@�`	WY%��7�����g����/O/)�� ��NFx)z
��k�x����࣍�+�����]c�;��a�DY�"àD7�Di�&>�cndNv�`gAB>�PE��t3�h���R�Aj�Q�K�c��Gj|���Id}��C��Be��;���
- ~�^���l�f��C)��Q)6*�m����P���S�'�D��mدn�3��8V�sų�Lmk�E��`��Q�N�p���C��O�?_oU�z__��:ˎ"�e���t��g�Tz�'v#O ��xς,��`����~o8���-�QKp<@+�_A8���e퍙�q-���E��8xR�Icx�EI�� �"�A	C��wh*&��p ;���1A�� �Da `*�ZjJA��G��Pl���7�������������+{d��f$�U��^��FW{/J�h��:hx�.l�)1I �6l���5H��0E"�>Ч)4	�sLt�vO�<�'��N��N_�Y�x����i����w�����/�m(J�4~/Z�+��m�	�V%�ؔ�fxGc��,ԋm��Љ�<���GN
��Jf>����N,%<0�T�}����96g`"tb����-�&�Y(�F=M0N�������/�1U׈϶aA;���%�M�����;΃ �E �M�l��-1�����`9Q ^1o��\�E���e���l��ݞ� x��q !_�b�6��<�+Daj�"QAY���g`Y���k#�<EY�d��;���&�[X����##�!����D��},ثN�\�O���_myZ������.Zl��q�n�m���IW{�,6���@�..7��M���a &�2�2�D|G�t��H��_oR����)�m��l�^�cS�t7N�}d��="b��zݦ�j���&9|㉉��@���vl@�����.�c\ɉ�� of_������AK��G0��m@� �����?
�-_#Hsc3�~�og�k��n�`��x]p��?�kI#(y��8�:�2�(M:�g,��̘!q<\7������>x6M'�,�����x)� StrL-�F#�#�����}�\8�ğ�Q��
!�1
xb��'F>�l��`m��(���f���I\j���b�8-2�.�d�ɰh�eޑ5�k4MM���uR��5]��I�����˳�o�f� ���+�{&D>,6NfzM/QSx�ᒉ�v��`rX�Ag���v��*"8q�b
�Hu����MV�������G������E�N��ͬ�W
�J@l� ƥ^�UA��u<D�q����:>J��dW^�F�tI����I�x�H���C�;���m��g�D��~�@~�e]4vxx�z���-ٺ&��U��}4.d�ʟa�+�Y�hb�W�_�5'���I b�$��k��2�#�B�: *Q���{s[N�ӿ޿���)���"2Ó?C�05ˇ��l^���z/b�29�Z!Pe����D�?�J<pTw�V4P��ڂ�~�)���|O�!��)@Z��>��N �Y!\U�ف3���_������ ��~�n���~x>ҩ%K���L�*Te=���%+�!@C��	�T���ↄ���\�p�V��Ȯ~�j��8�+&��q��� e��!��ј'˻�����Ym�H��^r,���=��XA���D����7�Cj�a $7Z�Qp�R;�@I�������ghs�4���-89#�M �1�WJ��O�O���?_�Sy�2P)MwQ�h�&|c�53�m1��� No����nJ)�u�"$J��h)<D^ɽ%���^�c���j�v9�$Vw�z�r�u��cZsN���I�bpG���f���{e�_k&jS�+Li
f���jp��p�T�x�mg�v4,1�FĬ��Ae�K`�x3�$vK�`���|k�+axk��h�0�I�����_������� \�y�� �� �A7�H�8j-C���sz��Ys��n�5����"�qfg��c��>� B(F5��Z�$6�tgmE��"���2����Y����@=}GT�.&-)`&Gqg��vR�Fh��k��M�?^	x�����ӟ�^BB��9#9gY�md ]�4��i�:;80��~�����}�1�x�3��)<�<]�⩱_?t.ێ�6����#rAЭ��|�3������zz�U��7̌	䢫+t$��8+�6ދ�L��5���<?C���-�8��7��-����*3��I۩Aɗ�-r��ԟ�F�]W`>������^٭��n���Z�O}�<��nV�>2Q��Urv���D�F\JV��	�!��O��'�{c�7�����pG�0RI:ب�Rf�Am4ιQ�*5�/���\<���"lD�}�����HO&R�e,>�d[�4�}zV� �[�M�6Z��m{z���� zJ"E�5��"�6FyAV��틁��CK�J�҈����t��&w���٧IU�Y*%JR�S��j����/	A�O�����z�Ie�@N�L$p��Rа	�N��.�"���(d�z��;x�~��;x���x> ����7&�UMj�M\�8���ǡ�t�J���t�,��Mc�]������u `����t�^_��c�x:�O]�)�eH�͙�od�ff��ǝ$��k#G�� ��k�6�+z]d�%i�����u�hIש��gs��$t=����?@[JhnX���i��]�ʢ�FN��e���v���N�mo�}?N��F�2�]ZS�#R�W���N�]�����Qa&s���w�3%��@������̧��|t���7���7�f�΍�(���o.t���:-�y��?�ڑ�4�;;�iY&z���/���ib:3J�E�2b�E��<�{�|�p�H�mSa4_��4s��^��r©�߯z͘,�y�N�����-�ݢ�?������߳UT{ܗ"BPC��̝9���Pȸ�8?�/Y�]�
˃��5UC�)�
ի	A����b�Z���l��d�������l��ǰ%2s��uLW��.˪���\����:%MY� E�h/�_��(��1��N�V	-S�*9>�m�w����*�=~>g�%���4d~�:������> E�	�o��f�W����H���,`<�t���Y�	�����Us)Q%�#����l#�W�����v#�B��ͅSu]Qi+8�kT�~E�qP��
�4�*����ָp���z���E�)
����wዓ�7<Ƭa�ձ������K��~�/��KZ,�!=M�0)m,?�b�e�P[R���P�`���$��Mؕ�OG]?;<SS`�)���W������g�"��g�QW�����'W�t���H%d�Q�o���g٦���k��t�l� �YD�>5�b����Y�����k�#Eq(+����J`qg{:`O��)���  qK7ZL��i}�KZU��8]FW��E�ۤ̕_��+���M-�i�L������8�Tsyz )�2��f�L��a�m�?��n�/�/����w��w8� ��0��q����3��~�d*�h�>|��%�6ؓ��p|��r�5�a�h��2.tE�[�D7�L	ba239v,�2-ʓ�,}�Їˑ1u#R<Sol0�s���$��@�=��l&�U�kq�c<�q+�	(s�܉�h'ϖZ��}�Bk�ː��i� �e�5���+�lf��N�5 ��y�FC�e�N�K�(�@�*uP�U��`]�S������(Uaoäfd2�
�`����X�ˊv*fv�6�7DX��":`�[�meK��Vs~j{�'��-�&�A0��Y��@�ŉ�~`��N�����e�	�p�6f~�{���AP�=;i��5���HY{���9�kD��&vUx��}����*�����7���pk<��ۛ��?�������*1��8��G�����U7�@�m 9���'�[[i׻[~����= ��	��{EL=G�K��9Zf�-���y2(�\��@�&�>F�(��`�U��jŔ���Q~��7Ͱ<���4O�;���!s9��' ���G.Bl�����~R�s� �D��w�7�$�]ebL�ie����`v`�A�P��CCW��[�P��~	���w���V[��b���go�D�s �>v����J�������t��I�wG:�x')()�'9L��r����yں]fIh3!Z��w|%f&.����>��%|2��ཫ����%�gpN/��J��Kg����}��8��	Td���:pf%lw�U����pɚ��ua�7~�xO�4X�����?���@� @�WN	��������Dqbh��)�@���|��x�=h��_�#Z��0i������Y�>�<��&�>����Ӝ�h9T���9:C�M0�'ܺ\�=�����"��d$�% z��S���ষu�;3,mwh��Q?��1a�Q��y����x�z�S���y���)"Ť�q_:ݣ`���p&�����f�2e-і�z/Q�e�Ǭ'π�jf��|��
7ܧgIA4lH���t�������2��d1�p���BG��C�v�̞`#��PTf��D����s���w]b8��鐫���e'w�ĭXW	����s�5��,��;�2:h�Yt`�x�A�*��&@����q�{��{�<��������Bj9�8�����!źc:5�K���)x��c;���Ҩ�4�w��[%��c��x2�?�"�43G��8)�)��.�}{�zp:q,dp:z�|�h���|���0ʝ�]3��L�Р��٪vI�9�+�S�57)��f�$��ܻ=}�n��������2J�@ft��gA����ږ
�lUk�]�Ѱ�d�@	8ێ4Iѕ�&�=�v�E���@h��@���]�O��=\�t
����Yڰ��@p���T������>�%��,
R�0Sdu��`���c�zU	�%G A,d�)]Ӻ�#�U�!'h<��G��Q٫M��)p�'���*f/��Y~R�?���
ZvH��p[V�
��Z�m��ӓ�rD�o��I�=,,�6���G��G �#}B����啈��E���M��|��OL �i��4l��蹏��.1%�J
�u����c��$�q
XJ:��3 ��tñ��9~����� ��Ԛ�TLk�Y&6�X�i	�o|�(c��u�Ee�ǃ��xx~�~��rD�s{_\C�n�ga619 1H$�:ڔ5��4a6���#hț4�hw{��Eh>� ��փ}̈J&��~Ai�( ��y����,�L��8bO�#^s��Nx��H<p,�&.ݬ��s\+���$F���`G�QR�D�X��B��� dу�����7�_od S�+�1����u�7�~�y��Uy��dd��yj�{u�C�"ܴ^�'�	���M����E�Gx��IE���ϗ�p:����o�����J	�t<i�cj5-���_���:
�tw��5����}Ɔ�9u�s� L0����x�Tz�t��� �,�Ѡ���6v&�Fj����\o�����L��}#�ΩL`jR�f�`��w9N�����nS��Nc�p߂��ڰ�ah��cg���e:�:|Ղ��P����2���gF�K���-� %
�>��|S`�|ı̗�qＤ����U*L�'�7Q:6l>/���H�����+���{qlJ�ǫ�:�,sW�Q��� ~�ER  �梯�/@�\j8Z�\�rU��st�FA�E'!	�1�W�HUb�}{ܗ��5�����p��JX�S�OR�s�/���^��,�ˉ�t�W�=�Ѳ}�:�֊6�n⁣�f��([U+w�������\<����?�j��������N��s ���l]30>g�A�jt(�����B�s ��p-%�Ү:Z�Q�h����pf�W�v��8�"æx kHjc��~�i���4��K}�(n�m�MN߰(�f$n82�	ʙ��[Z�u��N�H�b//?�����S�S�O���V��c��&C�$;|�]���u���q&�FqT %�#�UL�´�k{��%�P��{��Y�>��h������a:�X�dd���]D!t�\7И��CF&�,��#\��2���� �B0�u?9���#��B�ǝ�ҡ��l�G��T찘j���Mp�.M�ڟ��p���2��r�؏�2��,��?�b�/ϸoe�⸖�E�3�����k����#ؼ���5Gߟ^^��l�i�����z�Y�nX�&%$�$�����/H�A]͟�a6�"Xp!#��St5Y��,�Mn��XS9Ě�Ǖ�#K�Z;�$a)�h�!�;��� n@>���h��	+Oo�M�����d��U��~ěu�,S�j�����h�\�@�Ic_u)R�)L��SY��wܾN�hݟE�E?�L�4?���R��ޯ�=K �I���w��Rj���cA'+�L�q��nG���+��p�G���:2v�3e�WHg���Zaӕ(����s6��P.��Wy� t�S^�
����	4���;1�6@�@�J��޸����,���_%'���������z(��h�R%��N�m��ْ=N����~�b�^��/`9����j�0�Y�1'Vj��՞�o���&=@�|��lbb]5[���fM���p!��I>�o����H��l�UǅfdY:'����L$-�ϙ ��k���	Q��m��w�y$ ���e�����I�+?�o"��Xjutd�О�~���"��O-(,Vq����F˅��ư��6ݣh�|�X��0#�� 
��bydY�{ת@ə�=��4{t�Ffb��b��I�/v+�`�t�Ǯ��Ύ�Ȗ,"�'�X��?{�zԖ��G������=���R5k�r
�U�X{��h����nz��BK��|�W�`O�5L�%��n�M|�eY|��ԭ������^~|�V�Sf{��̝k(GI��%:�~��9<?=���Z���]��&ӈ�N ��'�p�� P�c|�̓����TY灘��y��{�"].�j�f�٠l]�OY�7TV���;�Y������߿���Eɑ�h��b99.����pI�Z�S��z���R ��Y鿧f~J����R��$W�n=��J�,V� � -}h��+@�PB��E�)CG��'NGg�+� 0�lx��d�>��h���+�]�y�g�wz��Z�E��-�Pz29���[�#qӉi
A����7� ~;�]�<�p��S�Z�o}|N�􍲄A�!p����1�
�t�2����wiB��K�"�7����^Xva'��偂m��I�q��`L<.2t;��k����n/_��~���:J��N�y���$߱q0��U8� ch�`�o_�^�i����O9���l��x�H[�w���a)֔�6�j��:�}|��p��\-���_@�5��gF͇l� �:���FԶ�����	�����O�i����A�����N�ɤ�=�6t�a���jM,��Zm\�}���=��;s����n@�{r���><&�$�6|�|z��o?��e���b�uMH�j������H��f;��_[|tO�݇m�7jܹHљg���Z�8x6�쫼<w�����N��h��a�]'��|�<�΢Ct���*O̘�懍�����Ʊ����\��52 ?@�����X������5��i<l 1r��~�w��Z�= ��7��i_�I�����S7$y'�Y����"�@L�����j��=�i���ގ�������M��15�E��O�f�����Y�#�E,�+��R�a�����g���Gv��h�R��<Y����ӑ��z=M���$�U���O��+ڔxڳ�P�����S�C뽏Q9�ٛ����Ł��0���t�*ˁY?Y��}����h\���w��3������(m�;��0�G%FKC��b@���wO�eo튮3����B33Nd���W*e<{�{ex�{2�Ԣ�M=��e�AŚ0�(��|f�wb4�i@���=��8����6�����[x}л�M��A�q8QP���x��g�7�g��s:8�R�=��4��in��.���'R$�`1��;j�'�Ssi���j�P�]�ڤ�X��!��3��d�)L�����s J�����H[~��/��xe��!���%*ir��%B���rYf���<N3�w��\>EP��Ԓc��O�r��������B�ēlE�^��o��?��<Ȳ�;߽����޻�{v�0�	 @�J�F*J���BE��(ǲ��U�V�*G���,��H�SJ�Ib�ab�%� � "�s3�}zfzz{��w��r�{_� ��TJ�0����������;��;Z^��\FD�4�i��Ȉ%��
z6��^ 8�Mc������T͟(�v��҄ G�͟�8e\@K�.bQ���p�3��(�{*B�6|���f$B̤g�
��x��Oh!j��F>
���s�E�Ԏ(�C^����/�� ���!������b���������Z��$���N(��#�TD�-��97�A&B�ᨎ�0iPP�9W�v6];cl���~�kq�2��6�ʋ�H˄���R|��>�)�gO�"f��=�͟(�F�O�d�Ʈ9Ʌ�U�,�V0^J�ـ��Go�kPI��
m�V��c�a����&�"���#A���@4���Yy��&���Q�������`(<D�z�Lf�M�8���4#!(�s�8`�@|7���۸+R$����3iu�<l�	���Xs8 S����B��|4< �V&*��:���9 ICKK0��N�w�'Py3�_;�(eړ��R�.# �1�ԋ$6�¸���hł���a'�	s�$+_�&q�	�Nd���*�Q�K�K�蹰
V��QS�!�b���cI�TJ����%��h�A:ɿ��TV畼Ďc̘�Lb�\T<c10�Z����#vj1�ť�7;HN1*>1�k�f*I�w69<�P)K�AJ)E�K��O�J�.�u%SuM$�|`�lȕ��U�*V�G���$�0�R�|>����5���/��Kb��+Y4@���g�sP1��:u`AzQ�POz���_��k��R�,iI��ؽZY������%Q�c⇁������K��ux�ˑ���P$P�ĸ2�j��7<X�)o;�I�5��Y`��2���yPud�%�y�,]0��A���-��	2�X��tm�6+�Z���CP�D�g�(�Ϊ7
e^�		��
���Eq�P�����,#��tZO�E��Y�w+�Zfc� �g��i=�S]�ae^�$�C��T�`W����:��>{�^y~LN�H�Dt�p=�=��2!o�E ÏU�Cփ�X����8S�b���ʕX�ؽ4��6%?/���׃F�i#o� ,��X�$�T8@r�=UMC�)i։ɏ9��L��+��e�o���{�̼�L<w[?����y���*ב4����P�{8�Y���&*ZKl��z�M�ڨ@m�
�A�Z�͜�Y�n�id�1�,���Ґ|P &�*aӘO��Yu��҅��2e��~Kw�-��D����i^�z4v���TV3��8�,}�tf�4S��D��%Eo�I��r�g��X7{���+�^��|���i��jLr`��RLP	4�ڝ䝁T^C"5zV�T0�ˀZ�rv�Z-��~�Ȯ����32�@dK�s�A�(WCX����T�&�.V�pj@J2I�(�Rf #hʺ��F�됪�4�� 
�
�(��G=�&O�#�{�^�#%��1�#���㾘����a8�k�&O���H:�!"y|��\"�=5��{��5g�2Je#e:z���3H�&�T+%F>�y�r�C��(L`���<h�*��d2@'��=�{\��%,�ì�(�Vz�TEs��uv�@��@���lv��S�L�x1	KȊf�8Do�0��ʡ&-�T�,���ǜ�2\�e�<W�fB�/��J
����؅�jV¥�,�Muѳ��ʹ��3oLM�m/d����n����8��!>h�|*t��@��R��:g��d��VC��t)�44�fQ�c��������[�*�oxo`d~��}�瘅�a.�b7v^�K��'/rv.E�cҰ�Z��6Q�Eڳq�%�*4M6.��f<,���T�~���&��S�^���&�Rx:]�0��$��A0U��&+(�Y72HJ�H�;k�IRqY��tr�G���UAK �$��4K���:4�A���iv��6���Ty>"�&�rᡨVEb���=�Ɔ�\?�n8̩֪0�l�Mw��	\�J.&�NQ:�˺�l�H���я��B̲�:\��|^��4L
\![�D�1@P|� ���O�ʈh�� g�l��sy*�m���ay=�(��I2!�)�	�z-wf����2{�{��П�n)U�QK'l�T���?��y�M#x���2l�M��f&��I��s`l����t{H�c�&�юL��(V`(���*�ݗLy-�ъ��`vx3��u��3���uj����P��"�ey;n����wu^��3��=B.V4u��lR-�Y!䉩���a����w����h�ϟ(��r$}
��t8�C�T��J���{�p/{CzA�>i�N��tH3���1cR���U�]�\\n8���soe�	���<���!�t򞶑U"Jq��D-����A�"*aւ�n�yUȚ�R�A�ʩ!�f:H�#��иh��sB��R���^��r�Y��܀H�hWH�?��0���$J��H��
�C/�%V��.���=T�1e>��jQ�G�,hv��i�ˌ��מ��:��NQ{�,���;�=G�U�O�~b�e"&<�24�}'�L��Y����I���*�&	\YH%m�rݲ@Ă�9i�#H���$ə��o�O)}��yƼ�yx3)(9{�|�T0�����
�^Y��/H�SREK�`3�"��N<-W#��:�H�ъ�i�(���O4j���>w�txS��"Ā��`�V���T�5
��� Lb`�3e*�-��=�[d�z0�@,��/��]X�zy�C��@*^TP�?�`���)1��CH�H$�)[\NE3�� �t���-��7�nf���ךV�b�jYn��n�,� ��$�"'ε�0�&�<'Z\)w�N��>)Di* �op0�-�|[C����QP�Ո�c��.Jn"��Aȁ&��v= ~���(��]�|��3�������%�\#�9�F+�2! 9����J�(���@[aH��z��^��Y1Y[���n)X�m^�'2),3�k��ƈA��.z��zfX$Vi�<e}��߀QwKa�@;\SAMU����c�YY������L]~H��>S�Ƭ�׊ѱx>e�j��p���ԩ�NSM�J����P|M�� Ú�M�a�r^���e����/eV��ȱ��V�y0H����n~�
*g��}&�TZ'd�˴ǩ�99�%��#���n��J�O}����'���DN�j_>� �!7	�Y��Ǉ��e�.���Z���8���ދ��tC��o�D*^�'�X*��Y����Ս�?$�e4xHP�����Y`#1��i��e�w+��t�sH*�L6*���[����l��RtRL'M-�P�9,Fhe]*��xIՁ���w�	��,˟�܏��G�$ ��Z%�h�d0DJ/̽<�ʹ]��^��Q�X�졔�*1>�6H:�)Z"�tQ>�K"0µ�4��ր��(P���g��<����L�{.(@^�x��DR�&h��J��2U�δ�O�s�j�·K�$���� 1GK>Ao����͍-�|qx5$V���223�T�Dd�N�T]G��d{�r��~�.�m�J��8>����vZ�ehLMC�g��*��s���5ԫ1�f���A��3��sĜq�3��Jy@!w�� �&w�|�jP�l����p^7Q���y.�Y
�Q�v�xKA+E?А�G��(PG�ǈ���u�u�r	�C�A1:�~(�s�א�'�W{oT�L%�2�J�����V��@sp�&в�<3��.,@�j��AF&�ة�,��	pٕm7��f������������Z��^~}%f㵰,��3Ϩa-u\&�����t^=����=y4�R֫�5D��|���BF���XW�(�¡2��-��D�!M��+���T-<�IX���4�8f4>����yq�9}S@�0ysrr�D@� H��x�g@U'j�B�V�+@�,l[+d���if�y���X�ϝIi%)�+(M�>-���:�4q'���5Nޛp��JFrs��B �0�.�MqRW��d�u�X ��d$!��Q���aX�&^ąS��FR��I��ߑ^�4^�e$L�*R�����X�k����I��J�M�Y�4��<�?el����|:�^�_:=�sDR#��9Ort��n(����x?6
��OK�A���aX�t�0X�N�+~J=%�iS1J&�bzO��ʡk�)�Z�`Ǯ-3�.(��p\��_��|�a�JǑS�m��A�Ӫ)Z`-��O�P�m]�Dk4Y1y��J�DN��4������d�JB
�K�Jj�S�9�b�$	�X�t�S���J}8�Ɗ����A�����:��F�����d�[$mR�oj���q���>a�O� %"����N�!\9�A�S)S��D�z���M��}�Iȋ����(@��ʊ�]X8�V�4�ݨ��`���[�.?�v�֒�P�`T}(B=o(���NoN�ߥ�v��r0�H[4�6t7QQ`�HYN2Fq2��LF��*��-�:���*<� _��z>ЍL'/�]P��,�o�uC�[�&Z��U��,���;99Q��bS�dha�âW���9�ؤ��f�Ȧ�)�>sy�]����3� UÜB�m/��+��Er�Gh�#�z�X���WgU:�%'g�`Q��O�WŔ��#0���nAh��\3�+-�u*�<�	�,��+����8����;Thځ�a�VH+��߼:[����5mN�Gyd�N���'�C#|��K����8��@�_��j�n������A�ؘu��UY�7���	A�S[Q^<c6N��2���|pZ<h'�Ci���b�b2`��;!_$&o��D�"��qtq�Tb(%���ZT�Z�
oN��F<VݩL��*	�T��E��]K��V1bO<	�(��<:��@΋eϛN��0�]�Y׿#v���,Jmyə#�L������o�V�0,b�3E���y�;���ƕK��v������U�zv)Q(%o/s�#��#!-���|J�d!73D�Tؽ��B=���� �
�6R$��L5�$���������b0�=�_�q���yEE,�5�C���㸤Z��>DVNh�� ��K�3e2�T�t�^�K�݇�̈́�LiM��=9�,��gXt��d$!KR���������|9'��e�J.�����]}����%
�Ū��E�x#x�HO�-G�N�h�+�e�L���$Ŋf�����UR��Ӧ�E�m㦺/��
^AQ�<��i���B�a<$�Qn��L�ՋA"���*�F� �,B٤ym]��D�tl�1)��B*�y����꬝� 1#����Q�?
Cg!�WڕX+6�0����Ո�"�G�\�LFz38m��I1g��
.$�^z�~�"�J�{�<�b=GF�)s��	��JF��
�t���HV>[�wY~.t���F9�S�����eڋbFǎT��9hT��<�)X��ʍ��"\���N��[�k����<����p�--��W�"�<φ�+��k2�r�Z-�V��3�*"!�X�CK@�u&{/+�y6~z��d ��z� ��S�g(0�~��*�P^od�8%i�X��ZJc��k.�^�+dP����-�:�8����rBի��!�s�I/)����z�d:��f��?:� �\�	X>W��	#kE�J/~ �{�"�� ?W�����"ĴNG�$�&"�Lu=�M�r� 7��wJx�y(��n��Oh����2����)�$pR+@��ADi9xK�p�!9�IU���"��3�&B�t�ن�hH��K9�eBi*�*�#
��O.4g���e*�l�fNբ�<m��ᥚ��cX-�1cyN���r�&�K�5����\A�=Y�̤WJ��N#��Fj[�V���<��4
+�	�@�rX�J܀j��@�ə�%IٌT���I5��O\D����nL�L���7~¥/踦w@*A<�Ր���R�;^�~����A�ډ�ؤŹiMCO�Zj��ev���3�d��4/�1��u�!�N�˲�kbхMI���p��E��� ƔN���v�=��>��l�5*z]���l,	�TB2�4����@Z��92���!�{���C��p�DN/��Y�p� Ŕ/�2�����܀P�#��,���W��%�t�HG�	JT�D�H�N����y�yg��v��\�W��I��#'�4)����l]���(�7&������ؑ� �Bұ��	��r����k�TQ�#/f������h�}^�� x`�UG�z�Pc��f!�I��q��b�Q6%} M}���(MY�M�H�W�Pʍ*��a�X�`҄cB��Pt0-Y�C.��v�H�#ȳ)��Ϫ�2m�G���Fz"�n�~�'�:*�M�dZy�N�R��R�2�X�
Bh5!���@�䤔L 0C��9�	L�RfR�#ܾ�[ (@׿)����'��3&�M���=��+2^�ݧ�s3R4�/<
ˢ�@����T1<�����*ު�)׻�0hD�@��@97N��C��x����?Q�\Ԟ�dU�И�÷��ἥmD��&�ML�Jr�wd�
�+-�K�.R6�T�mF� ��>�A�J;��s؝rY��r%	#�S8M�2�F�"Z��a�������M�{�邃c�!��ű4�p�}<̠�@Dڍ�VE����ˡ�!ip�C�JF&�Ϲ�Q\�܃4d�@��J�����A��Rn��w�5� �,KY �va�y�簲��av�W�&�̃�h�9W��O'�(�	��u����dh*��;�.�0�KM�Q��!��44�;��ҁYU:8��Ɵ ��bL��� A�9���2�6g��\�kA��� Z�:�pU�5��G��~H�&��i!�+�&��51�8�.-%���ϟ��2�GV� <��*/�O=g 7�[1	�6�7.qSj�G"�jYR@n2�԰�e}M����DQ�OH���y�$Y����Of���A�0h�S��"+�F0���ac�y=��2X3N�{�.�

�Vl9*�d��r��0P�i$1y�b������JIǠ�����#O�QpN���>��X�� _O��!.��p�D\2!�� b�u`5J��^s��dQ� �b
=�&�T�Tq��'*_w��Ha$�R�)?�"����Da��YQ�7�a �����hu���R�NL��8�Ls��iHh��@�����7�Sl ���&o��6��� ��j${x*�5H�T]Tgd۽��i�WK�ҕ
`��BC�����T#�)�]�]�#!�-�RWP�f3�u�)��� T8ŋN�!@��@�
���1�P�c�r�����j����I��Nji��h�A_[�M2_5t��`bTs��1�@�7��`�ƽ`�!ѯ&�wg��`�J�m���Oc�k���	ub{^�ȫ���4��jb ��s��H#.�$6'u!���!qg�6����3�>\�������B���yg���=G(ɒp�*��U�J��*�Pԕ+������R�쭅�8�u����0`���jBW5v�*S��#/ϊ�d�ex�k{�#�R/=�!{|���m���0�	�{l�w�f�N4_�|ߜ��6��Gj�yӫ>D����B�6�y��aƺq��t� #?�}��4'6>A����ҧ�YM'�U���&R�L�w�\��'�KNS#��(sJ�{*o�`�N%�R6Σ ��8�Dd-z�4�=��H+��q x��˴d�!�1Wi)s��D�*K�"�D��5z�#l	��yd����@>�d�B�`o�A�8�A��@�9�t1w�2�V���S-;�N�骔�8xV(�i��mz�QX�0��0W���_6xM�1�He�L��U�3��(}�
Ʌ�Y`�7M0B�	��.i�7�af֕��84�6����碖�p �$�����t"혋4-!tZ�(j�AZ��Z/�!4�)��O�X�-p�J��u���3��ޑ�6�\}��3$Z�	�NW��i>hy6Sٶ|Ы-o��ϣ���QI���9�bD��2ٚ���6���m����/��*>��d�΋��y�1�q���e��������).W�w`k�f���r�Մ��������1s�U�B��R�S�y4 ���D� 9l1�ؐ�+�2��L�"�#��.��e�RvO���t����J�s|x҈9e 4�v&�`��VL� ;w?s�)]�
٘��Uju�w�!L��0�B9]��r�{�I�%�x#!R�F9��rjY��� �Cr�^�m�c!�� .��L��Vb�wӖj6<�Pj��v����bE�G��k�Íd^��HJ��r̋� n���Te��U��$���d*"2�.�Y�dB4jѵ���KI��0��Y�,k�7�H:���� RY m^�QĜ4�����	h ږ�o �g���'�7]
�
�ٸ^��2��H���<%��Z�T7���W����c֐E(�}6��H�oIAxv�/ޓBr�ͥ�$��Ʉ-�?�]��	�J��%*I`�;��H <:?*;3��ks][����!ɩw���8��H�T�|1��u��^�h�x
��4�4���U��j�'(F�7�}R�S��\ew��@W`�3����r9`�O/�.5C�"�&yt�_tMH�YH�<B�ۦK�x8�J�|�M��.�k���A�.�T~\U��CmC�im>3�I�d*%|����E��_�����m��ʳZԖ��?��yA斿� � iʨ�ZCb� &��hs`,>g<�ܛ��t!LxY("&��U����BM�,�-�T(�@��0B�8tE����y<i��84ʹ}���ѩ�"�@��tA2*���kZ�s��b4JK�Jv��� ��*!Wtx�im9�m�ֽ.bg@Ɩ�Ir-tV���@_�S�D�2�����|�U(b>5�>�cL%�����E{"N�3(��U6O�0�HE�"�sWgp8eOb:��"m%���h��B[�**�}G�轮	�0'/�2�n��C�.�2�y��:�'cy0v��P=����?�5���;��bl;�Љu�5D�}�ݏ� �<7��4�7@`�U$/.��,��z��N��^o�C��:��P����2E��A����ȥ����,�BR!����h��D�o���ᡩ��EuJڏ9侎ܻ[7�m
�������a�11��>?�׀3�bh��!Oq��D�THg�xU�@$��,6]H��7���~¨S���)_�J&���K
����ڛA"5#_�}	' RK�����2��D��ἦK
4;a^�*� :����4,j°q���$�,4�p��5�D��Q"�6��Q��8=�(��Fʌc~��r)����%5����7�)W&�(]#�ܬ�N�!�4P١j��N�!pN#g�#x�hv�I��pD��N�f�� ��<�I8�����6H�e=���I(�K%��������3ћ��?�����ϧ�S'�W.f^S
��L8	��B�X^8�彆�#s��u��D���"'�0O�dr���\��I�H�E���W
6�$S;�%���]��T�Q��.˾ EHF�W>�]ח�K�T$PK��U?f�NNO�0�w���D�JZ�@k����wEå��z5��щ9UZK��M�ȳ/�=k�Ѐ� rC%�`�����#�萮;��e;�Ao#hъ\)��y4`��i��)����᮵E�,�y�d ��� :h[��{��O���l8���8Pv��\�M�r/�`��O�����w��{���Z�+%��7�):�dt�p���,D�����t$���6�ͳ�!S�51�	�T���k�}z�e
�5?�v_�zU���.z�d��ә^k%C�=.�zU�YD�U
V��+DJA�����( 9���U*h�Q�W^(J	u6kLXx!�;D\��OȷFJm̐��(�'J�h����
:��8)��"H�)����X�����B.%g�J��U�b���ա�/����].���cd�Q��>/�ey��tq�O�"���<�7e0�V�BnX	L�,F����AZ���.�@���	46��I;:1 �@�B "Q���`]��N�����N>0��E�%�4��X��O['eeJ�K�|W��H�{�\�,k�'�4*�|Xvo��$]a�H�VMB�g�VS�'6@��`�M֥�iåZ�&�x���ɥϰ����q1~�����w=H�=��)���<�eut�(��9�
0��,��O�.�J@�%�� ^���K�YoB�w�tQ*�Uh0��1R�I=��Fͼmր#7�id݉
V61��O�'��y���g��SF��t���zk�s��ZAT�����<]�\6e#GQ����2J&�(�U�!��F5�!:hJ�l�I�O��\���H2��zc����c�	*/�w6�â���Y9�|f�n[��f����V����D��h�ф*5W�L��"2n����k��C�!���4�*4A�ݮ�2���@Ra
��3����8����P��S&�o?��TY�6�Ϻ=��y�I�"�P�}:e8+{ս�2��+6�[�$ߓ� a�;m�^K<�Riќ�[L�!9�
��w��ށw�\��2�Tݍ����K	��ҍ�Ȁ��l�TI#��'Û./����lñ��h3��VEHkя�Ò�'��ei��}2A��)��� Дm{���#�[y���x��P�Ť.-�� �CzɃ9�$�֛��d����9{���Py��9#4��*=|�U�!�8���l?M�m��[S1&�B��şVX+dކ�y�娄g�6����&U��\������V>s�s1��eJMu�NjUC�,&%��i��9�P�e^Y���+��I9�tc ^��?�1�k��wX�c	5K�!����tjd�	��R�����d-�bac�I�<p�$Ay��H�`�l֩�=�w���� o���-�!��C��.Ŏ�`��g��{ �F��K��	�Ų�@}?'�p��5�>pL:��-×���*�����6�D�?�,�V�@Eg}޵���,�7��Lq�#�ӥuUBZ5���$�b�1U��y�<L- *J2��戼M9��K��A�,�}�@m��U�
��9�ԬFr�)�� �:��. �b�UK�<Q��^:�UpN�5�@¼Dn�9��SaV#��&�k�?���%�k�6��3=-�G��Kt�S��0���b��@[���gz�z�hID��s/�#;?K) �.����8%\�!�(G:����>�M����8�H%���c�:�i�����gP�;cR�FW�H3a�^�U�_�LMG#��,g�;+�{[3�zqצ�m�WH�"4���!����!|���X����r��U�����F8a�%�6z\�j�Hġ0KH	HOc����$p��k���(��OV�}��t`�,��$����������˦�����y���̉�Bۅ��Rx����+ c����$M%�f������52�,�H8��q��Q��5Y��<��]7���V*s��������W:��s�j�4_#A��M�&�I�'�iK��CW��t�����L?���2�ى��`�~1�$����S��	N��H��.K{(�F7Q�3M�T��p�^-�s�BY�ajA�8���)Ӕ���{���Rr��}`rjb�R��s�R�R���%�z- S	�U���d#��V���ai�PԼ�T�H��J�`�Q��VD鋅h���'��HXe��,��x��a��d���D��rz2�L���yx���g66ozZ���Q���M��.�B1��٨�B>O68=w�����*Q��N��L����8Bg`��q���9���S�G�ـ��{�X[��/G�?��d��(j��D����q8���\:�=���x�F��3|qP�/�q�?t<:&��|y]�Ƃ�,D�	G:��Y�����cN�_T���^���V�������لLR>�B'����HQj��hfW�/t�w�L$%V��2��Е�ƻP�	`ŭ�*U� ?D�C��շY��j+;3��)V�nD��Ԥ�_R�cZ�Lv=ݼ7-�2��x�:���6.
�F���7N6�c�Ɓ�y��'񪌫�҃!�QS#���R�R��,�6@�W���VF�aA�u�&�O��｀�H�)�n!=�����eDZ��6U�[JO24����r뽑������aw�ٓ%�HE5�{?��)Ss��c�˛�V&8b�&؊�Q��th�~H�YVx?a,�9qB15wɋ��6�{!^+lG���T��a�����K��Ճ#���o�!�i��=����q���֚�u��Ox��,.�6����a%p`� V��E8	��J�h�Gu3f��k]X��2K}�UR֜P�,��r��ߩ
o�^<C�X<ǋ�ay~�J��-� �Q �̀��3+�C��F��	���0�k�0{4j���Y%˃F�Jg����j޺���y0h��VPP���w����(	2:��ˈ79+X۹��В��$C`Q��6H�B�ϡ�Y��'E���T�C��R�7Q R�v�o���Eȶ��&����`M�Y.�(N��-�Q��b~"5�:H�� Q�y
��8,�Q]�ЫE�	EH17�c��D oo��H��܎�RU���Q��i�q�k6� ��q�u��XK1$�݋G%�y���ϢeN�	�x�]\���&4C	SI{<�Q��L�7�,�c��)�����8��ۅ�{��6,�'�큏�:D��	�3q�N^}�տ�w���S���,�D�x���30fxO�c.G��-l�D_u�fE9I�<,S��,��qB���L���%0�$��3�ॹס�Z��xdJ^bE�2�$.��a�-�C�N�t>����<��x�-h�FY��S�,F� �*�C����F���7���W�N$�f\\ɘ�~��X.[e�4�� ���fZ.�h�\?J#�֖+5?9�`h���,V܍4l�q*��4|����Q��h�h�<��+lx�#��$��K��L%���3����F�<q4D �:c#2�0�n��dH����Cג����Eߘ�%*��Q%i ܈iRK'��3{Q+Y���F��TR�����!�_�G�I:���[ǭ��N��-�vuJ��10�6e	pg*f��!�| Y�PI�}��%xesP)���>]oI�x$��]ޏ�N�L�ϻ\��L��P���gZ`�X�'�%)���`��T�����|k	�8x�{n~䗡u�c��F�Y�q�ر!���OG�υ�c���qO���
[ag�t:��a� u��\�0��������\���J]S����Lô3*�v��zol�͋��l�׉�s��d^"��=����c��8�o5��&x��t�Q�A-�����)���^o�x��*����Pm�B�y5媣��~��{}RiE�;�b�Qa�^&�OhϾ�x�����7� )�YoWT�����*U �k������׆�zZ�l�o�p����QJU���}�V����4e������,��c#��Se��\�>���i�9��!A��
�� U�=c�y����*d��ZV/���NA���mطw�?�tI	l��&۷p�Gx?�R6�}�g1LM/B�9-�F|�m\�>�9�㽽��Gb@���y6,�J�\݆��}К���;�h�0��b��3&|�=��C���A�`c���)XZX�٥%�lw0GY����s���ü.��Μ=���)�h�c<�\eh�Z,%G��|MT��95�W/rd���y�]w�GϠ��a�C�I�-(Ee�F��4�\���z��Y����4>��ol�,����%����uvJ�k�����7��߾K����kB���Ӈ[o�	N�x���Cn�kk�}¹�af�	[[[@m>չ�<�2��kvff��accv�=�z���ռ*�+0���JoԁA6n�,����;]�Yy�4;�s�v&���0��:�אָ������'���;3}���y�����w�.��ד���~����9�kfZ3�����m z�ӭ�C�kW���\�����_�9\(�1�qQ�;b�/^=�ߟ�ٹ��N����`�-���1|�XZ��"���<-�m��	�ʱ����Q���Sp�] ��k�4���gcq��E�+���&@gϹ�>�������iX���0���iY�s������`~��Cy~��}h������`��^��Kp���p��]P�]�3_���ŋ�a
-����u2���:�B�t�8��(�:�,�Y�+��{5�N�Ih?��x?�檰��gϞ�����=^\�����x��Y4,�|��M����WV�W^���h.��E�355��-�%8y�L-Ǩ���8�v�<�t$w@�:��� �K�h�h��ht�5��`��l	��C=ܥKW`��c��K�F���O�����Ϡ��}]`V��J�Ԟ����44�(5�P)E��mh���^�� v�¸��C�*h�HBqq�q�A��z)��񎧅�&'$a���ՃP[�1a2��xf1R	ȍd�;R��1Fu4��^[=˕<��h9d�Ҵ��0�/�Ti��ǭ.��Q�7�p�?�܄�C#��,�ȥ����@?�ZU!"�����8��N����h�l��:v��n����h4�h B�kL�0%��ka�=Yu�i�[�.��Z߹�M�~��cm��7��~*i�T���F��.u��۷�������6��배���j��?��%4ѻ�����'[WÛ2�
�zʍ*Dׯ������-�h�=\��Z���X��, ^`�֐B�Ao��nua��:L�M������鴹"��Z� ��:�ٹ3G��ҽP-�`�vN�uH����0�bp��)���EU�������kb4P��$�qcR_� ��&,UC���5|��b!�L͢�;�	թ��{��=hBS�:z�7��><�2B�zV⢨Q�a��=T����{@�ʆ����J�2n�ZCp����C|��<��µaO�kx�����h���9�Ѓ��\�	0J(����c���
>9���^�R�:Ԧn��G�`�}�\=hr�<�0�B{�}\&�DOw�`���mÁ[n"�3S)x��)%��Z��F�sK��c��:n��2ohLD���9���f-��0"ᵳZ3z�2FG�阫�)�$��*�_������X�����M�1R[�C)�8�Pӆ�䂫MF��H��k��Fb�,F/3M����(X�'4H�O�N�� J�az��Ğ^�X��c+t�6<�7��$�B���ϧ���ɗŴ������ �L|ԥ=h�R�2{�8�r�C�F4���ҍ��bb�����/�ö4���u8D������+��z�a*��?�9���㯁�ps������L3zצً1?�ʮ5� �IQD���m���nDeH�[��q
�#��[Qܜ��Dm�t�0l���b&�9̎bax!�>�fӎm���"�y:�Jy�;K+{��_\V&!���^^�+o9�T��MC
�+2��=�r!a��+u�5�㨛�v l�A@ �Z4�/�T�h<k��z�dDZR�e�~�P�x�xޣ4��ln���^�{xFh�|��Q)ե���d��A΁�� �=h�kw0�af>� �JD�f�D�ч���P9>J����҈F|��Nm�n�(	 �ƨ�*=	k�����{O|cd�v="x/\�����VW0 �����2�� B7���F0@�v�0���[���E轢9e���Z�ǀ�|܂\�ӝn��1,�EG�i,4��n#��z�:��4���"%*L�i]�JV���6b�4=�@%42u,.i��ô٨�y��`|��ϥ�F#�:^� S������QU*JӘ�A'�h���%�,��R�|؃ '�"�m@�4�#�Ц����@]7��Jko�&nbLY�0ŭ��q���}��3�2�_�U=��~���Jƛ�&�z]�1�a�zMΓ@�� �xy�0_~�t��pP4:tWO�ǔ8�()�-4�T�b�OF���x��� O��g�Q[�ϐ"�<N�e��"��y0$Q��Ȝ�KM���0�n,J�x��2;%�y�0���7�d%������z�#D�\ 	z�c3��b|�ۇ��4�E	gg9n�Ѓ�\_��)�,k�`����=�q��B��1�u��C�� -٤Ri�Ψ�d ]?�k�����MDu�C����j3�U�""�u�%)�4c��1T���s���-��Ѥ��j�a�:�A�B�/�[�w:pi{�i�^�&M��5�|�=�@���`��"�v����7S��`�P��+W��B^v����  ����4��/i�.�Y���o��fC� [��G�De޳87�p�("�{�&f]�ĥ^�$�8�_��.D���'i�*��G���S�c����.\�ف?��p��͹�p�q
<��,�F��ַ71������<zb� Q�G%f��L�$�I#��e	*mll���a;48��!Gj-|~x���A��*�6���G��������F��tޮ�;�@�M����n`�h(ʣ6ۂ���V��Y��|�%��Wavv.]���]�W;;8z�4�c́��a �Jꘖ4�}�j-�u	���j�����̙��|�@���;��{����PG�2UY X(M\F����Q���n�� W�?��>�	3�Ȕ�B�i2;����������5�%g���p3쟛�~��-8u�ط�Z�^��UZ�;�.���������5NaH�5&�@�(�'�a����#�!#����S��~o�&��!��<�S�9���L����`�Rܸ��'�r1��q%� @BޣPT̒,˥)���,Ѣ��6��ns�5Xǔ���e衱�֧�M��U���ř���J�o���W�!�Qy#RS.�W-�a��L��`*�:cI�B��Ӷ�)�4�2R�f�*�*\S;hH�ZBU�Fg3h�ޮ�;�@�Z-xe��F�@  �����\�a@��Kd����;8�߄��S�uƃ�\2�(�S羍�3������x\\%\���Ø�y�َcrL��{�oU!�P8�rڰz�
\:�]X���p���ȋd�UeYE�����hpKn�Q����Ua��.�)1t�=u	��F���M3���G���u|�`�e=�v�k�&��� ���vJ�Fpn�,WM(�	��s�>m�hc�9��	�@�Z��Н�*���C઎�m�
е��_��䙫P��a��@�T�!RZP��PX'WO����F.4�ĹIu�'Q�R�ԍn��i��Ɗb.Ա�
 FB�}d`��������K3�)��!��	���HҀf>`TG��z��^�[h�:����1 �A�<�Pi��Vd�����0)�2(E��&��	Tj.7Q5�>޻ J�ѕk�`Ou
F�!�]�w���Cتdp��� �F�4���^C�#c�'��Ha���aBUr��nhx�v[��F�V_�׻̞�X����x�q�M-�W�c�ڄ2��}�<׶ס�k�o�sY.������PP���s4ô�
�Fo�y�J>L48����}�#���o��r0S���p���hcj,Gpla.�x��q�TBh�w�jMC=W=\���T4�w�vo�a�T��@��Tқ"��H��Yn,B:2n}!�V�hĺB�"� 4�e��J�L{��a��`D��	���x�vpC���@R��BӼ�����T��t9J�=��T!|�R�#�Ai��a1�9u8���E��>pC�����A_� ��h�1���I ��^�f��:�vÕy8qm�G�%���@P�p�7��u��^�	�	mh8�!��H��Eh�5	1�9TbHL͈	F��F()���]�w���M<���ԣ[��E>�0�UR�	R'jYh(F&��T�❸���y����BА1����q�x��,�m3{���Ey(�����h\G������?�����M\�	4j��������z6��� ;�1Sc�ݻh�hؚ!,.�{o�淇����p��"܈���c���˗�B{v��_z�U��p��w�,��d��1�f	2'�>�\��"�6�D0�Q�Yx_�PΑpr����7ie�5�jj������55����e���a��`�����U8we��&4�`�^��r�� p�����QN�Z�h���@�D*1����D�pR�!+�A��[P��������1U(���1�$��Z�A���ȫ�VO�7N?��a�<�������B���T�J��d�����[��zշ�~mQ��NP4h��w���n/Cx���ۆY�a�Gz%�U�������͑e{��7�S��Å�/��ۏ�{q��[��gn��~�:�0���3��L�Zp��"l��]8��)������Mh� 1� �=�2)���~��T�|��^)D�y������p��~�����f����o�����֨ϔp*�>��spi�4\9w��.A{vN�v0Uف*��'N��{�$ ��K�$Eǀ��b�NT��|��-�G1L]��z�~x�mwq����z�3-.`�c��q��/��<\�4���k��7��QT�\�!�q#2�T�#�x`I���C{��ܲL�D�ռ7p��%���<��0�Da��A�1×�#j�l�=?|�fسo?|��/��Bia�1��C�Y`�M[�"�9��a񈜭B
��q":�:g��r��v���w��@D@� �q� �nE�,�(��q �d���$hC���s�%M��6EK��@}��o�������5��ōF�f���Z^f�(\����!|�����>�'p�����p�Z�U)2�i�uJ�N�D30�3r�7�6`~a�-\ن����]��w�_��ǹ��Ҙ���n|�^�����u8������߄Ǿ{
*�aii�o�{#���V�!� U?�	"�xJ����Nw<4/m���G��w�g^|��'�=J�;��ԑCp�M70���ڀ#S+py�<q�[����0�Ѐ�L���V��p�#E�ԇ�H_�iCH�Z�i?#�psA���{�}7��k=x��'��v����p�v����ˇ�����;��~	����|���p�}�8���#X�� vd���[�O�jW�ڨ֥�ׇuD���
��H�K)z�n÷��G"��֭ݝ*<¹�
�p�Hm�*�y���>jW�����_Z�㛫�lÏ?�cp����KO<s�J4��+����lcz�������p�$��۝�Ͼv����~����+���*��sMx��N���e��a�\�L�v�~�0�<znnn������������<�ї�V��{��0?�糥��hX�^����(yWc�Џ5J�������������7VOB4��n�y��N]��ן��U�=.i��ř4���q ���N
?q�C��c���N]���N_Z�j�6����z��ՠ}kԪ��=���v�~����d�:�l�b�E	�i65߅�����35�a�i26n�:F0�`zԼx~���G��|��W�o<O�e���w��م�����:�β��W�U�<x���̏���Om\Jk�7�CD�>�uX�\?5��χ*B4z��Tl��^�l�%t|��Uȸy�"�@�-�4M�$�ѻ�7���w���١�e�2_���U,�t�9;��t�*RkNA$"u)_���\(٫����G�pc���0;�8z�������_�7֕�J��A�U*W���?��v�����?O\<���/M�LM���h������> Z��Wp������^� ���/����G����������򮝇���^��������Z����N|����`�0�G/���F�⇷��l�j�~$s!J�O������T"(�]�H������M���Oë׮�������C?�/jP#&�]N|�����V���������#���ν����y~����k0=[�n�C6���9�k�،Q_
�K���3��aa���V��;��]�Ƴ�\�Y9����G���������ǹg�y��q+�쭷�뷿;�OO-��T�}����n�1%l�1T9?^[�|�x�֊/M���(�?�n� k`֡���ޮ�;�@P��^�����A�pS�L{6EcT���H"�^����f��@���U�yz|���K���ٙ=�'������qܐ�թ������'j��߼z��w�s?l�!\�����p�N�)F��)�#�������#����^��[n�3׮���.~�����y��\{�ۢ�������o4��觲ͦ��!l�҇��n0�=�a,-�$����'�؋�r��ZML�޷xV���ĕk�z��|�}�~��u�A̡��>�췟���^�'��||�T_�E46��<s�4��2�jhi���jhw��ѽK����h��0��{�%���v����7��?;q��?����y�s�<��|���ӗN����������6��AxS���Y��Z���&)�:��z�0R�6�X¬�0w,)�dPB3�ښ���u*�F�;�@����ћ1��RnN~��1{`�|G��=�E���^JUS ���H%�
���}�b������~�c?�Kh~��Ӯc��\��v���F�_n�/�t�8���\�l3����[F�b5}4�(y��0P}�Y4t3��n����}��w�{������q�<~�����˿S*�>��协���yׂy��K���Ollqw$��4A�q���}��7�|R�c�+0H���{~�ÿz�����O}��_�~�����V�D5���;��B-�C=a��0RϿ��~x���G��g�Ϧ6��{� t<ld�Qo��/��'���'����������8s��V����Z�,�Nc4 13�R"\��Q���P&}���F�FiX�����Rv�_E����ӃH�#/zk%�8�U�Q�ƥ"�6��M�v�eQſG���{��}7©����G�C�����q���_}���;���j� ����w��9�zFZ�C�����3�G���>�����m�o�͵�����C?r��ޟ���ޗ�����j��T_�Q���knX����߫��,w; 7b���KU�-�qc�Fh�Q������Ax����|���y�C��������x�e}���!Xj��;g�c7�E�{��'7��B(�vm�T5�JJl�*�.��^9�؞�}_3��7:�}�}8'�M��׾��k��8����"LQ�k�]"3M�I���
H�A!F��v*����E!Y�"2�y�T6~��o��i Rn���������)d��E�c�6C�Qy�Ml�8��	��c3a�rF����_�7|��F���/����*S?�8�n\>
�W_b,���@W:���p�n�k�`9F�ߘ��Z�Ǟ���V�:���)��{�� �z�2�~�)�	��bQ�Q��M���{4�C�i�r���~��\^��@��ɧ���A:���x��&�7����
��C�3A�Sa��*�
�߬Ee�.h C��]�n�+��/>��?;!���B�:7.��{1�������H�C�����?�N���SŻ�<�J��$Un�d�c ��z�#D�����4��A$��tg~���̊<?���k�Ȟ C�
Ɣ5|�#��<��0LN�E�/�l��!Z�)88��s������!��B�7�ҟ�

RP�tXgta�
,�p��M-�a��?������?�����{�Qb���H�E�ǁ�����{ob+׀vѲ�=�h��𞰠^>�V���ݹ$M�v�V�{B���p j�$��cQk4M�M�Z@)2^B������������>�Z��f8\C��Jw��S��0�B��8U�'�6T��p"���t�S�Q�8'��i�(�+��_��u�xa8H���KpB��ץ\�LOS�<mI�Vu:	�����4%2������Dz��U�2���<V!..�r�T�|���_"�i�(�-��c�Pa�:�E�v�hz˷���]konA�����:.ք,���H\F�q�@�.��;ޣy���~������.���4x3���0qi8�#4��{V8b�ދ�&LR��Iz��z�eh��<�@��-�_�Zm~�>����MO��ŵ���N�V�,�RZ����xZWYF&�>��,
���e��U�|M��)����Ἢg�U�{d�@ ��2Ì�ˤ�ۗi欤�e9@��4E�z�]_.��V�3���+1��3�ݳo��h�~�S���]7���O���a���	�"''f9W�sa܁�ބlSzGH�1Ղa2<:�!���+��+n:J�q�	�W�B�Ӄx�� e)�U�[f�%�*�Y��q�3.j�:�Z����>�$п�Q+��^>w�r��A��w`}{?#�f+j<#�APn���td ($�cj���J��������O�:EE6�T�x+���K�)_Nc��o�����-�.<�?��1F6jR^o��2U�v�=��6�9���%�J1�5��P�8����xg ���J�b�:��H/q�WkN!5�=�bb�c�Y�3�"���)!5˕��������[ݘ'N�A����a��\�v	s�.D8�,y��#cn)��>5��fv�1GG���o�|�|ѿ���<�������N��h��٧�
�F���12�+��d|K%�H��E[���0��ˏ�h�������Ͼ�������^o��ݘ>��� -M���hf3�Oiw�e޾�g���i6���p�(~�%����{V��@9�A�߃1�R;*�A���t�sU�\��
Z��5�^�@�!�U�|F�ʊ�˒}XeLlD;�ᵔ��Ĥ��&���q k�m��pppn	^~��O4�����w��������m~n�� rp��y��y	ҊcBИgS3;��}qn�+e�����:�_Z�o��>�o�����'��}:{⅃�y�=��h���:���ׇ�]�.C��3p�MI{4�b�tI)v�5��JS�V��?��o⏞�����|��Sxjq�^��66�`�׆�L����WA�=H)&��^�-�߰�m�ոt��/>���迕���g�8u�������"��{�cX	XU�U�(% �*���C�����q�\(�<��3. �߾���{f��-M���2����g��˲L9�̃z:��ưtƕ�:��ά��=�Jp`q��ԓ�f��3�3�珽�:0��?��w�����?��񙓧�!�������4"�|� ���l��m�����I��ݷ�Y~����S���ѣw��f���߈���o��{�o������M٬��.�T���B��Q��=�D���:�f%�55��nf���_��7�����ov�������+W��#?�����\���W��.��Z09���Dn�dPEt�Hf�.:aV��N���~��W�{�̙3�u���7�h\��d��_��/�k͇��l�ڋpn�5X�DkS�����+?+"=uB�	��T�d���H��*�	W!D�(ʷ��4��\1�E��i o�����ГrY26N�@J���&ci,!oJs>H��Y��;}��NA����9x�ŧ��������g>w���\��W?o�>���s��fX*���`���kp�o�y<Ǥ>� uK�o��{|���Zց&��=�P�0�������c�~���W��x��?;��O~���g>W{�����~�#�p��ix�����Nc�Ro�j{�`��kퟄZD��Z�e�*u��6�x�ԙv~�}G��K��0��3g���������ϸ7�'kk�m���?����ܯ�u�{)������I�j%p�R���,C�B)^�@-���	�VX���~n�]�?�����>�	ȮmA���u�����u�O<��<�s��d|�3�	���z��V�������\����9�gV[�K�c]�����P�,'0�4���R���i�u�iaVN� 8� >ҿ|��H�=GJ�ZG�1��k�-H ˙)��
YN^���D�:.A�V�f��$���w_��������s������7�s7,�m]i��J��^�����?���Z���?���O�܉��|�2l�7`g*�EG-�#A����	d佷��Cs���!|���K��$\~��9~Ӎ�x�����ȿ�ꣿ��^2�8?_��2\	��_z��[���������7!�SO}.W�C���Mq#�#<o�Pu(�KMS�љJ؍��N�F�������k��B�y��;�Η��Ǘ�?����R|c�A��Ш���^~������_���7���
|�[_��^�с ��� �V���:`�r�ӽ���lFҌtp��I�g_z~��A��ظ�X�������|�s���G���|��F2U�.��?x�����v��ʃ�\Z�7�Å�9��)��Z�y�x�,�1��y����.�OQ��{��$�pA1f@0�Nd�1����2�_�!#����l��#�����,]X������I�hH�a�Ŝ�O^��ڻ�9������L�����RH[���dPl�"� @�H�������'��@$8�a;�٢���Lm�C{����}��7g�U�M�A� 
A����pf��n�{�Y��}��ۯ�>F[��ul�~�D1�ߌ[��:��kƝ�Q�\��'�o��A?��џ��t�[[�q���΅خ�b�Y�?�8����u갺k��e����.�0���3��އx텗���=���\~�R����yz����{�:��xǞ����֟���~����~���F��u��lJ��vBe���˚H'�&ڌ���!�F8����� ����W_�
.?w�z�&�2���7OGߤ��n��á9.�;:-�ia�����Ǹv�:�O�C���b�z1B�T|�����L8�0����%x�b�u�i3��W^CҤ0�� Ս�%,F�}��F��5�ЋYj �`�L^K��;�n������s�6y4}��J����u_�~#u�D�4^����:��71�;� �9%��=D�����+�?�,�2O+ )m��.N��H�}G"+��v����i�����fϬ-�?���G��/����m=<��:_�.�_[9j��,��_��Ut;1~q�-ܼs�������f^��"���#E�>���*s�8���p�����O���K��j�s�^��vo��n�7}
j��5]��6�Y��S��8\����hr�V�,x�@c�*�;���@���܈O�����o���᳟���{���B��ؽ�_Z(̳l޹�5������:w�Hr],�t�|�y��@`�^�ݏi��>�_���L�Q��q�k%�b��ʝ��\��Z�[o�D�RF��\d��9o��ZL�;��u���|����5��{�3┹D�:�1��}����hj24�px
��T�7�����Ah��F�U�O�(�(p͚�c�/��0Y��U�����5YB�s���H����9�	�=z���J��B��ş\~c{�b�A�cZDs�
��Ǎ����!ų�}��h,G�[�`wdq�Z<�iWd�1V�z���N^�7�=qH�m������Օ+����_��k��N�`{f�T�e�6�t-��8��8nb�T6k�Ў��d�����E�]zA7�:T`'�4fy&f�eM2G�xГ/��0���>ĝ�/�����xy~�b�>N�Z莻�я���9h=@�vP[_C|���w�G�C�/�3����cFhFE�A5�aS��c';�۟}e�
y��1�uT�[7�a�y��s�M��Y]���;�?��GǷqpr��t����gJ�Y������ǩ- O�c��Q"S [F���T�xRM�f�$���Ii=k��dEY>�c|B���@�.��O�\{���T����b�%.ԶM���GS�f~��L�ϚQ�\�v�&�2�[��]��W��WV��Q����g�����N�G�m8���0�E���آ�pM�ذȗ���O���ř�=���WZtQ-�ws=�/��|��K������.c�4���@��S�c�N+�����i��WPow1>��¤��1���3�	ǢI���2�'��,��~����g��s/V6���gQ���ݽ6Z�%�pB�|��4����%��*�'�4䤧$�}I���v;�.� ڬkZ����M�qVC"���y�����Z�_�x	{�g����<�A�s(�0Zi`;��KvN�p3� l݌tMf�R�c"�dͿ�����3���\���D�^j|m�b/�I����4\�Dw}�� �Hf�lH\R׮�[3O*$b�@G"�QY�.FR��ze�;�m|�����xyi���6�8�����:�3���d(��%4��q�>�3�9aL���������L;l�Z��m(�W�\�&��N�Ůy���5��_�jTB���)�h�h]�i1�ѣ�;#o�Â/E�R�8;�g%MMĹҝ����HF��>k^91�>�{C4F�x󬁅�X�ɣFS-O�I;{t�<�^�>�Yן�	}v�1����|��Pc�F��G�	$����$��+�_��R��4>%
{��#^�͓����oa��@�%��>�5:_d��udqWk��:>D�K��xX� JX�F��gQ^AQ���F��y1�Yy3��Hᚌ�>���n���SN�O�`�����9�"�:u�R��$I��D`�^�j͇���j��O��/��m�M��L��+a�����n���{Q�@q�M�FR����"h��=D��(e	����4D�K�0A
Y�R����B�JS]Ā��9��GIK�Ki�Z(c(�?���(|�0g�ꎝr\(Rra����`�HE2mb��:q����, �/�c���|�K�|��+IcS���5�vs�[��U�{r��\a�3댈���`���ą�Q(��K��kX�ɢg ����W��ha�Dcp��R�6�2�h��dh�&ᜄ���rY�1���4[����`�À���q�1t(\6��)8��Kfǂ����ޟx�ҹ钓��ׄ�?�Os��Q�IR��"F�����9�'�{F�O���b��*IH+�@�Mi'�!O��y�W?�,��:��R�۳�x�+>�
�[�[�UÓ��ﲬuuf�U��)ݜ/�aR��}�8�Ї�����^�;��kk�8m�F�����1!U6�&�h���ɉ5�Nb�b�a8k������w� /TA:]Y���2S*�Ъq�{`�igP�)?��& v$1y,�$�E�ጏ�	��V����P�眇㥰fy~cC��|�a'�����2�}�%��2��)-Lw�T�qthR�f����_Ӈb���}��{Gs$�4��ө�w�MS�=a�Si X�j8�~$�x�
q�T攰��wE0�X��.Wafp�7�@2n�n갑��S| urm.��5��������|eWU�ݲ�U.�N�a�få� �S���m�sa��A=<�@�	��o\�QX&/��$��5)�� D�a�b%ER�jb�)������\MʢM��]Ь�a�_��oz7B�g}LG+�;K؅S��ܱl��9�$�fDC4�="������MZ�p�n��;}�j\��d����+��{�(y��F?I<�2>z�@[��@ss{��� �`r��>����4��0Z����z���ߒ;�Id;r	&_(�$��E�D����1xz��ɔ��ܘµyu�'U��jDt�1(����H?G�xgd�z�� ��92[�ص�ٱ��,5(�i\3��Dc,�k�����Y��kʬ�M[�d��.��*B�F�R�ȵ����*++�N�F�%�}�<�@�R6yi�C:��1{��$-k{�W�w�UV�2��7Y��惬��7��d��L]��.�����!����:�/QK��X�(GK0g>MR~�M����p6D��x�$5�'@l��lj��S�G-lOMl�0�3;v��p���}��O��e��ylՍ��ݵ-3���-`}$����B��Cl�����Ȯ�6�0�k2n+(D����~?��{�c�ѯ��x�07��Jr0E��7��d,JWt}^`]�O�����rw�r�&���ԭ}D�H�'�__<��{Ϥ�N��@J�qKhl��,��G'-�O{�b�*O���u&\����y�i�����~-,a���I=�J�-�^�rW9�kE�y4;����$��F��,���K�:KK��-m����&�p�{ӿ�K�r\�?84���Q����gǮS1m̶�@���YF�;3ag����q�`��ĺk��?����d�-L�����<�&���y1,ᝲh}a_������<f�#t�g�^�����Y+��7:V��e(�_�aXN�&��=.$��`D X���I3�j�8$�7��xrB��cVfq�gl������ � *���ȱA��Nb7�%��>�.�y|���l��?�	=�J�p������n�o�PL��i�25O�
M$��,�.!�b!8Yi]��5��%/`�=7��v.g;��%('�
�	I�Ÿ����ovzYxV큑I�Ju7�c�ʎ<O�����i}��O�X����s`^���S�����"6�(y*��_���Q<��%[M��v����#�
<�j�Rp�:��I��Ӽ�+j�.����;y_!��h�bU��P(�g*���y�2�B;+���E�d2��$63A:$��X��w�!ęR�R	�ٹ����R��J���-]�H��}?��a��9� �й��z!�w���k6\T�u�    IEND�B`�PK   א�Xw�'<�  �  /   images/48eecc1e-62ec-410c-a9f3-e9ce63fb3255.png�YeTг�%�nda	�E��kI��^b%��K�������.i�F:������9g�3�a��7w��U��qipQPP�d4�I�?����w�U��8.
n((H��0�o��?%5\V��l��p�F����9ٻYY�Xs9��f�Ҡ��~T�����:21�B����l�1*�(WH���bZQ#�,Q�Q���C��T��DA������I��׃q�t�}��1X���PRj$�km@���1qd�j9r��YG��]�~�Y���WX�z=[��5ҵ�� �G�2Ǧ&��PI�c ��p2���*t���7F���3�7!���X �R�Q�n���aI�2v�̩���A����99��}�w�ܦ;9�l>`�E��8�������Yz��a��O��W�q��O����:3(a�{4
�u��Wᵋ&̪���F<{�j��kr���[���mUY��KR�x�P?�%�^T�H�m�^����?�`�D���Fm��H�w�⡂s��&L��B;�Ґ��oԒc�MR\���������![����Mb�'�o^u��O0��'� LP7���9X{^�=��c��m�(SL�clv=���п�-o�I���QRּXI�)��A2�v�����?�jj��G"�Z�\.gۻ�)F}{��J��� RΥ��b�zL(�;1.��>	���Y����^��cD>�A"��f����Sz]w�m��a����8cAeE�ʽ��8�+0��Q�
A��*2�<Q�b0Rz8�$5�9ˣ�U����t��/a���F�$���>��ăU��VD��aa�}>	v��
E��幫������m%���iW�:��	o=�{m��ڜ��X�z��T(�^�xPG1�36WA�h^����aqly���RY�?�����Q�1�LFv/(]��|=��jg��X��\V#s1π��ļ�*�D�]v�o:��K�<h�^�Ә��nO�[��
�X���Ɏ4pc�8K�S�p�[���*�>�;$	j#C�0�'�,I��3gIi��F�U�E�k]wS/c]p�ܜn�:P��8�cn�0�_�ު�T�1�Sa���)ۻG8�,:�e�PQ�ƛ�Pd�:q����B����U{`u�g�`�Oq>29�h�6����%��9�4HO���7�(�_%)#U'b�GY�O�:�9�W�ܥ�7��,�]	��S
�2l��|��z���]���^��^��Xß3����f>�(M�r�|�5�K�&`�|�v���Vz�Ԫ�^m�y^�
��U;�&�����&�U�S�'jϧd��=�ڔřQEh�%�Zfp*q�TTg�`͂��K.]��ǭQ����1���䦭|��&�Y�o�HĈ2�$�ѽ�嘅*�<MJI89���9�ֿˏ�X��͗5�������Q���Pl����}Fn����Y�w����雅&�|*�V��ee\������#`K�7���di�/@�H�ᶗc����� �2f�qp vug��>�V��u$�*H����Қɕ�����n]��5��*�Lb@*~�Q�Ah� V��9`�j{��
��@N<4���p��*0�r�y�J۰�1� �Ef�pZ�4d�f�5�L��F/�V�@�z�.�SLeC1a�H�ڍ�B�������~���ݠ|A�� L�Tx'l*��GG�]�!�3}��+Ղ�[����<�s�<w��4�-F���"w�J�\\�!����Js��x�;�t��e����O^�皈����w�f�d��/8β	{ύ�IXh<Aͧ]�"��[՘��Y��n�?�c��ގ'�����$Q���k�u��J'z�5����'\�/��}M��[!����@��my�w�v,�d8��t���zrH!J��/�8�9ɯ�smdN��<وD�a+E��x�0���8f�����c_����n:c}��4�``b�z�
���b�D�P���L���@j�R��k��q-�O[:?�)��+�MD)����tG�X㾕�D�]��2ڟ�*)�Z�dxy۾���(v4==�,���o[�T���QbE`TfD1�Lfm�p��8��/{;��Ze�u�s4~���ī�������uO��cno��o�OX˙,p"�m~��496lNRU-��go�`�[�G�j��3�az�|1��6 1����t��M�+���s���Sh��5�?O�~'�v!L�n�p|�c���@��ޠԟ�g��P��7�aY��]��"�P���[f_���7H�\'�2�y������pM��d�v��NKѾ���<��$��6E��#�|o�t�7������v�?�N�򕋑)������(��̑�{�K��V������1bM~$�ل�*A+6=�͑u���6@gN�ԑ!��g�"����Nh��b�4��r�5#P�>���g�4�ӛ�q�ַ/B�z�a`o�6<J��*�mt��"6����N���ö_��|q��/g�1��M��l���5f�n�Vs14X�,,�l��F·����S��})�v������Ppy�X�:�N�E����%��&/�i�l�����؝>�~��{�=W]㉞a;2S�1x�G�y�M��|���U6�-�H���]��ơ4<+v4�ae�1e'Z8�Ύ����~ȿ�3M6&��t���$k��
K{tg�X�l��o�!Fd��Ż$	6丌iho��7�����cO�P����J %炏�{ 6��Z����dSk�W�qO|�:U�̇�	�߹N:g<�JO�g�e߁�{��Jݦ��UBD�'������T�������䆘,aI*է���^��Cn�<� Oj��;Қ���bU���/����WE�t�M[aam�����޴QY�v�ɧ��8|~�L��6kI�&�|��݄��ز
�[����4�l�۸��9/o���Q&�ox,bOK!:�ՔzX<c��IB`	����Ѧk�q�����N�|�Ƕ�]|����4�����jx�=���G�݇��_ϐHU'���j|��Sdot>n��Zg7Wl�룳@��n��`.wR�vA�gwRs�m���
�E���~��2UDMjH�2:x�Cӵ����*�9���E����dɐC�S�K,66d�!�1���Xp�qS�#��8����1!^�,�̞�)��+�0GX�`Do��[�w�k���*�Ŀ�v�����o��*��7�R�-���v��gj��e��#Q!~��?yxW����}�����&��֪����CA�U�%O��F���-�E��a���K��Ծi�q�uS�f���G�h>�*�1i���
C��L��&����zz��O�+�/�]}p��m<<�XfRX��'j)QL�3��	������:^tű�q�*�PQ�I�0^B��l"pp@P���,��-Y�죷$�7+���Î���a��SЉ�vb\7���a�#f�.N���e�G��L]��$7��Z�m���2���Y����Xf��^��2�hT���(��O�)�%ԊL��W>,
��&��dm�{�ew�>��� ��e������ǅ�m�qF����{f:���l2�$�vf"kb�C�`&;`%�����"��:��c
by��C��g�����´<�]��~2�o{ ]�/�(u��<*��~ �e5��D��6�ng��}�~�p�D� ��+Z��N�f�>b�F(qGg*շ���s�$n��5/�������Z� ����҉�ٜ¥2���1�E�����pW��,��ߠ���n���[�p�Mx>��f���xd���$P�a�q��Y��{�#���M����oi@LnU�U�b)��՘��_lm��q00tX�z��JU�6��[c8��\r�U}{�y6�awp�P�Q9���eCe�F
xD K&Q�'}!TϦg�����2��o������ٚT�u�G��ő��/"�2�5�F�e2�,Ww4b��e��k-K��7,�BM-s5�/�&d�Kͧ7�\��c���ù��v
�޺�iI�.��Z3��E-'���_����'ٔU���*�� 3�{��!�
��w�L��X��
Ņ�!8xO>]�ԛ@��_o�=<0���%������P�ph�H[��]k�9�:'X��r��l(N�J�l���AQ�Jd�qjQ���YT	�M>��>V'Ts?ܫ�\T�s�H�Ǻ��"vʛ) ibF,�1}�NR ��c�}I�L�C�Z�P��P�MR-?=�qP ʕM��*P�����}5��TG'�9�J��ᐒ��ˢq}V��6܇蓜�C�aT&5��2��Ut���-�#�8�m�؛�)
�|zMP^ݤ�;�+���ZI}�������)�u�,�3{��{uE���6^���p����d'�	n�X�e�~Y�GT�b4y���y��4�@D�e�6b��%����r[hH��7�����4J�67�D� �;���� 
�G�xBm��z�o����8�vp�s^���U�"���!}�%KL��c)d��YЄ�����6�.?G9|��0� ���f���ޜ���u)��ڤ��G,U�:n�T��@4Ck�.��b��#��D
��EA�s�s%(��B6G�s��o�x$�!�!�*eO)Y��N�٧`⛉(>��W�F ��A����M��G�f�+�J��ƥl)~~�g��J2C	vh�n�?0���Y�Z�㢾r��?�5]Ei)�0`1{����u3��O�xF;|xE3��a�w�t�7)!"�R��`x[P�^�]������"2�v��Vd�"���=����i���'<��MQ�Lh�11��Hb8fc�3D�j�,UM��1$�f #�t��1��>��P��|�oZp�����|����Z��@&����\^����j����F��a�+N��aq��%jm�Pt���p,��@���)�)�ʳ��戟6���I�s[s"�E�t=쁮7�{��X_����1������O��I#���k�W!�^���
#�j�c&�Qq�I�ʳP}��C3e~�dZ��E���}LH��	�΃��O`�j��*�MA�߿��"�r�I�CzS�~Y6M�
�7�J����n�*�Y""�3�L��K;�V�(����M{+����)Z�%�Jy�ȣ����T�M��{�ai3�Ǵ"今K�^@����V��(�����/�-@�5���5�a���CD&#�'Zkn��Ԓ�jf�z(�E���o�wH��=�RJ^��������V�9�h�7^Znt7�"/����F�6�o)WlH�*���Vx�3���%>l�W_�@Y��$8N���e�Sw21E52��g]/v�	hy����c$�9{�r-4�7���[zw��:7��7/�c��,e=9L���Eyx���{��ũY�H|h/�
��0]f�(��|�PX;�����zU���w�%�}<IZ��d��0�;�me�z� ��/��̈�2,�n�3����ǟ�ا��:}�E��a��1��*���������,*���cĦ�ȋ�ʩ3������S�T_�l�p=*�UjY�J<SI���p��yZ�5�����W{|�\	✡�o��i����>6�����a�W{��UB�H�C�i�� 0�Eg҆�rԼtf�h�V3	���P ��?����0�D�#V%��0����~@���R���ՠ��b�v����w-|���Y�l�D�@i;� �C�;W�T��c-��H�&Aެ���6[�f*��}�Tj�7/K�S��~������yI@�<�^*�y3���8ա�^�r�\s�w�z�I���&��T2�ۓ����7�����2��`�=^�X�&a'�^��𼓻S�p��/�n��v���ˠT��H�qi��#�l�ŝ��ܰ8��X.gr]i\����E�~��z|���	����l}
N�	����Ki����V���u�hV���^�wv�	����~sCM���
cb.�����"���(����n�ޢ2Ck��l0��5��Bt*n-I��CFR��9�i`���C���,f@��'�C�̲= ��į1�$���Aπ�(�y`��OJdD�q���zO�b�Ot���,��=�-��EO�޹1��qa)�򞑧�)w���ٍI1O�d�##����rcǑy�u$�6����)퍭:F�5��и�|�=��8�դ�^�~�К�!%�IZ�$ �ز�W���52��sm��fx�#.MKw<�ǓwT66����0E\�k2w�r�$%{�p�B|������b�>9��i�nI��j]�K�}0ߍU���[�yTήzM=�y='�� `�ӕI	u`�r*�[�R�I����ߟ|)@Eirx��4 �я39¡ۻ6�.((2�;Ȣ�3kO_~��i�:��e��u<��u��b1���+��V�$�hUh�gB%�B��ߙ��ǧ�6�}4$Y�9j{1*��m��c�@���&��,��u˱K(tqbV(�6��������Υ|���]r��[Wtaq��Z�d��ی� ��9�U��N��,����uy��-���ȸ�����E@5_?b��A��'��eun����}��;� M%�9��k���z�:�h+�̟�w+�-��t]vh��UN}�X�f��P����Xn��UZ�M/�F��fn���9G8Y��PЋK�]�G�oւ~�8;e,�=�>�Y-����3�l�/Q��Y��I0K�mL8�ķ��W�{��^��L�A��&���u��k�:V�k�@	s��2�-�hm�rO�Zܺ�q1�=��`�HkL������=�D￫�#nk��f�7?�ͤ�|���/��6Z ��g�y�1
�ތ���J�_����u���Υe�T�Q|x~�ՙvm���})����H������qڑ,(r��Y�Q�R�>�lrϋ`Sg�}��Z���+���o���ׯ9B��V��2;|=�|���m����0��7��V��d~��]�)��V�˥�0��/4�e�BF�� 3o���C�~��'&�����������=Oѹ�_���<�h�xh9w���A/ٿ�ޚȟ��7�)���ş��G}P(qt-���uB9#�-3i"V_c�"�S�V��%�C�)�����J�V쀵Þ�Є2�If��Qt��]Hn|0��e��r�c��#���5I�L�����Tn�)[�o��]Ჲ��f�X��)b�3q��T�#~��[�*T~�1���=n)7R������ë->�R3>5��(�*S%m�?PK   �C]Y�i�4�6 �6 /   images/67f527dc-1a08-402e-85e7-42fb10b753e8.png @⿉PNG

   IHDR  R     N]   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��_�y��3�F#�XZ`&�1�Ǳm�`�rw�¶�m�m�[�-�m�$�3۲3h����}�s��H���i�d?{�s��{���;��J����g�������g^�q ��i�����T�)�jr�%$'�����i�M�>�/���d����X~��l´n~P3����Ɖ���JI���ƉMҕ�$�^�����;����,�&�]/z��Gi��<E��=��d���t�Ӵ\���/bs�sl��M(�K�>f�qa\\�U<n�yބ�����LDK	*olb�~���F�,�L�¼T��{��耺x}���� aP��
�t,ϸįA�M!1ʅ_�7J�N/l�����>�S����
�TG��3C�������7s@:3;mɳ�ʃ0������� U��'/J������8��e������ ���\�S*���x��q���Ó�n�y3�{��ů�:��<�Ɩ������Ƴ0܅&4	��zM��,(7����u����zַ��������.N���\��1�5Ԙw�������^����bp[��eH�7�y�R7�_���3�����ʂ�p��^���+��Տ+�NG��4��
�#��4Y��N4�Ӳ����$ɃWG\?�y�F�1�GI���ɒ�8?�������.��f�3�Q�yrZ���c��?�E1r{���4>�3���o�2�u��.v�������ۉ�}50z��úT¿_��?h?�Q&<��`. :�)��;o�hW��z�|q�ď��.)U�	�Ly��:"8�����	�JJ�	e #;�R$�(/)�[V�h ����^	 ������k�ϫi���'���=�b�����N�;]]1\�Q��M�=&�_h1|�"KY�n\I4�u��12���y��E�_/��b3WN�x����p.(ŝ�+	����H�ǐ�8�
j���3���Y8��p�_���/$� ]�T`��,|q��0��RހR�s%H��.�5Hm�Lx���R2�z3624n##S689c���62%��dKV�S��BI�Sަ��B�$�de6�u����� bBR�*��$6�u������*��W��.^DU�?ys�m0�}V�&d�%�$)}���$�KH���i�#C6:>j�ӓ��f�&lrb�&��mfb*��,�Cd����)�zᬜ��˷܂|K�Ȱ�$��(��	�?z��~�Y��49I��C��(a����#]J��笋W�U9''[RRЧ'ޅ{��+�[H?�;���2��}�D��;9�nR�q��N���ljrʜ����W�$�.����{���|tu>�-�v��?FW����ZF|�%��n/���/.���Q ����BH���b�k.��@���d��05X���W�A���Aow���lHgfC㙝':�`�;����_�GOXCK��u��̸�'�f�0u�� e0���\�E��2�Fn�s� 4P���jXj-��ns�Ge�s �)���ML�v M5$)���	���ɲ4�)=-=�r�m��dZFz� .��r�����RR�'٦&�m``�:աtu�XO_�utu��un|!��� ;����	 ��F���]��I ��)�i�
�''T���Wn� �8_\j�*�����-�ZM	''�t����N)�DKKKS�
/y�}�
���(�7�
�¦�T�}�}�I�Y���񛟟�Nޜ`<�(����wPn"���V������������ϔ����*�tǏ��ͽ��{���H�3����+��2NMQ�w���>��gܣ���d�yY�Y~�j����ā��?w/���v��,n0*)JSJj���_1
Ӓ2����_g
� �x�Sݒ&���6Bޓt�sLO˒��x;�?����Ġ����5�W�����a�R��P�FFE+l��<���5����S��m���y���;o�C�6:0b��RdgN�$�g�>W����}�/��P����"�QZ]c$�qq��Z��5���������Ժw�{�F���O�嚐0��8��qK�[ZZdK�*�jq���>//��垙��
N��%���*[4���qkhn�v�i]S����Ɣ�f9$�	|���fu��t�5�O�"��q���(Y�'�[��q����(��쌀zV��p�^cH����D/2��#�����PB�����"v���/�*��$��Osn|���_��|���k��������ziNsqE�cc!�!��z/Z�;fN�����M\�*|��Ge���p�%G�xR&�6
;�\X&~��Y��ΞK��Oa�HZ L�E�1-�F��:}u^0HW�j�3����w�HL�t$
?3Ŏ���F�{�z&:n�D2<)Q�(>HJg�z�2��YiIV��v��ͶjY�M��ŸP������"3���l怔�Oͦ�pӎ�ﰇ��em�Ö��o��'F� �TЀ��Q��*|�i�،��e<���C�pG�c|�	�{zF�S`q�p�7��w ,��g&";�$�+��OZYI�-�(���+.*�L�����62<h#C644d���6<4";�D���f99y��Q�YX\b	�X�E�==V������cc����[&�T�&��?�wX%P6��nb���*Wm(��ƃCtO!b��HT�s�*�:�@RvAPn(��I�:�(��G��!2�_Λq����/JcHS��8���G �Lz�߂D{2��韻W�)�ʟ����Yo�ĭ�r^�P��R�'n.�'NG0���U��T�1�Ɩ���}{��w�J��r�.#MF�&
	��[W�z�����|M���䑂� ?I�Z��]?"���+��#ez�H�b<z�:5)?�(�x�N�X�����8��]��2P&���C�l�r$�]�a�������Wm�ӄ�f������!c���5��tJK�nm]c���L�M�dڐ
tX�� �ЧDdӳjlp��� 
�f����u����N%�Ƅ�/�n����N�9Y�-��)��ğ����M��ht��ɑ~��N�5��m�z��E�VT���y��1;z䐵45��萇�H/+�4M�)Sx&�'��68(�\�_�d�U-[fe���SPh	i��P;�ĩS���c�Ŗ���zrr��4Yq���H�8��\0H�H���❎�#YqBY�_h����:�P��S��(����FaQn|��w�e&x�x8
�C���� E��^�>=ʄ���9�>���)�B�;��i����rO}�X�����@���߫�MN���j&���G�
h������ׂ�|qa�|0w�������r��A��z ��.z�s:٨��4�Ri�xS�R�$��*�i,e�����M�R��C>����B��hfE����*��Ŵ�LN�1!��7::�:�̜l5����ڑ$��tE;" ���$�nm�ܴd��~�g������Ci�w�^��3�����m3ǑN��fӭ�mľ��;R�f��o��6�7,pJ��H����h�������앃	7������FD�8]FI0s���mtEg�
 u0FDIԳӣ��4����M�X^F�mQ/�~�
+��U��g5g�Xݹ����#�>E�}����R+()�����j�I6! ��;h�]v��i�nq�)���z�:�X\i=�V��iu��6>�bc�Ӗ.ш�iX@���������� b� ���4o���@QA/��7��~� E�,#�ظW`]�_� �|	��(.�7j��!���s�I��#AR Ґ> ���ӈuw�"
��p�]|�q�Љ���6�}Ϸ�t�	HG�=�ܣ[�?&N-&��o��<��Dy��qnv0��]~�����4�wVy�髕��cÒ*�9z�)�]�3\��Ԝ^��&Y����1�V�W/S����ۥ����vB�ffv���(�z��32{W* ��J���:K��_��mǵ[����J" ��&�%Ўr�n?fHQL�$�Y}ː}��]vT@��Sd#SI6�G���b� Rב0�Q�M�ȳBTh4
7�
���dA��CBP8��U�8�r�����T�7F�Gu*�OM�͌C%XOXqn�mX]m[֯��$kkj�Z�h��z�N[.uӆ��z�r+,ȷ$Q��24���Ҩ ���˚����ѣVs��%��/*)������V�6dM�}���o9����]d�#��@t�a��E�9"�;/"�#���H��&*/o~���|G0�O?��!��/��k��^˸�8?|�WHen�H�<5��{�Ȅ�9�*-�)|��E�
�*�S��w�s���.����2�����tD���5�7�9�ÿ���ؼV>���0I�e(������� Z̑�o��q��D_�Ťhv��G�N�e�d��ۜ:$D�P�b��P�iQ�S���q&�j�t��;�Vo�l���TAɩi�NY��(���������173�;[l������}����k#�C��!I~�f���Mh���D��
W�iK����ʓ;HS�JmB�:�3��C�e*�	��{i"@:�o)t*��r�&.
?6��=j�&�h T�u������@��V�iUʴ��t[�Ԩ�[\��6�]n���j�ؑ�mbt�V,[aWn�l�W���_h)(�!>Uh��8!~7r���7.Q�G��ٚZ;z�@مe��Yb5�v��I}A���mB�6�z9Q�=r^�t<_�(��9���"S�:��Jx?����)��� �!�ȣ��@�Ռ�'�n�Ǉ`���aŠF�u����{�[�v_��i$
s�������|�x�,��&�%Wfh@��e�,�@&�=\lT>EW~���U!A�4^��2z�oC�����|\�vWq(_q8�zYL�C��F����Y�'���Gu��;5�m��B[0H�SE�fVV��1�&$ ʧ	h�����N���au�Ҙ(Pe�9���R%�A�*$%jV`>l9�I69�m��'�7دK�����ӮÅV�<z��4��I���?����z��عzkW���%�L@Mx#�����"8,D�n���{��Px�?���;�����8���A�Q8�}*�������D´�%�R���$?�VVU�-�N���sv��=�&�۶l�o��6nؤJ/�$���p`Ct�Y`�\�`�RW�Qќ�l+)*���|�s��z����ہ9?7G�l������蘾I���:��2��+eH�n��y��(���t�Mޣ������=/zC������p��U-�h\��aݝ�;L���������1�C�Cz��������i��4��?ᅐB8s�F����+i�&x�����2�ԏ���P��,+ǹ��˨��װ����Vf����;9�O�����c Tn~U���Ƈl|���Ӭ� �r��򳒭8?]��Q���3Rf--yFW�\��g�Zz��K,�GY$	�o�g'�n�r2�,S\niI�D�|�HO��L����w��plP�4q��m-bl��믱l"MzmB�[�(�`���㏸Y��
%׶�}��k�tqT3)�6�=��8T�g��1j�0!1��x��7�`B�_h �C��!D��B��b��Ux�v� > q5���e�S�x��M��Kl�
�ގ&;vp���������+�Zn~�%�f8�1�>Q ��|�e��{z��8���s��9MXww��۷���;`c"���Vۤ8�_9bgη[N�bK�.t�419]A����q�z�����A^��K� ��RP���B�`�̽<��y��A�{7�a��]n�A?�]�V�~�_q�x"P�?>�;�{��/H�;��ЅH����3�ޑ��}���x�S�HKp�\q��������I��ϯe^�-�N���#�u�Y��\��W��Us_G�MOي�EV^�m��j��6�(3���@��y��A����a�a���纺�����F!"KIK�Q���y��$�uL8 �Ԏ?i��V�x�uN��Y�� 3�N�{ɖW����G��0[�4�p�戶ɀj����ۯ?�9R�N�����X�<G*ԑ�0�'¹I��T�T	|˜H��.$#wS�^p�
�����  ��9��'�����p�
H����l��+�����f'�)U��o�ծ��z�ǈb.zȢP��R�	W����z� �%�@�<� FeedZ~N��I����CVX�I5��ڤ�!3/�^�D��a����s U~<� �~�'�a�>\��~����LÝ���~2��{�*?@He��y��w���%��wԏ�1���t�7��7z���S�i��E�x�K�x�u��L�D��Ǩ�h�t����U���� %\ʒ`]ݯ�Ra����Є��kX_��]�l����U
�G��P���Ϟ�(���	3�fff�6>hi	S&���l�
��A��ku�rie����̖���m��fZ��ˢ�t[T�gUe�.�-�(�����YW���L3><h}ݝ�8�|жS\gOW��U���*�{�)?;Æz:�zǭ��[�2E�6�QyG�(���P��|�DH_ԧ��᪪��s������?�?�`]�����8��{_��(<��L��i��Aa��zf�'����@5�ʭ9u�&GF��n�k���Rs�٥�����5
߼��*��+d(߇��(f�#VqI�]{�U�m�F�٩Q۸~�U-.�����t��Ihj+|@�#�g�`�Y�ѹ�)�+V���Q���[�P>�.5�o�P9�>#;���Gܱ�߂w�Ͽ��xl��P/��=u��aG��BK��/z��H�w�J��"�5U����'V�ͪ���|Y��e�D���2{"�w����v6!E9Шs��w��NK�����9�~�ߋ�.i���:Qyб�����s(+l(�_�?+��t�n2Kh��0i-�g���U�؝�\c7l� �=Ab{�-�,����I�x?;f�鉶jI�ݰm�m[��dڊEE�q�b[\(.6a�R�G,O�e��p����YVҔ�[^eU��r�Xw[NN�%�Y�ÝbPJ�>�\�.�b ��kx��~�MU��`Ċ�J�H)SrV��D�"�|�q��i�R��Lç���Z �-�+� Ń+���e�qu�7z���oSR����D�Ӽ�ӆ�"�����4UlR�e+��EŶ�"W��k��k|���W_g��x�����)��&�1�ڐy��c��m�>�&rU��i��uMqUAAi�]}퍶~�&��햗�fw�p���fXOC�͎X��%2�Y��AʃR!��P[�<��HY�8��˺�0*;���M���/O�J�JxjhtRX�Hu@���7!����I��(�Yʛ宊G�`nn�d�vphJ�گ:���� �p�`7b�OW����<�Fn>� H�P��9��y���YJˀI�N�xO�Q��0#�lu�'nR�üL�_��O@�,�|��7pQ�j���^���1v']��	�w�/�,ӆȏ��+�s�Gl�.���:׏r�E��$HY��MY��oTgɢ��qKNp��looU�S�v�[��
�FtZ�l�*�A�KMϕ�!�N�Xna�-]���
�����8d�����!yIS��4'1i�VQVlW�^a�]��*JJ,]���&G'}�#�
8�1���Wi�e�K�T�&/#�k~��_��*�IL�8%�Lx�����5Y�A�J��S$���#�c�oR��3jdpL��[�F��%4b���V\������~�c���%R�������Sԛ� 1���Ш�)�b�$%E�j����To�E�v�&�-.S.�j�yV��B��@�9�˻�s���s �T�Y�QXRn7l�L����U��rٙ�>�퐸5)Bx8���ݐ�@K*v�P
P�X�t�N����w�0�C�Y3�b�>�%�Ϲ������bآ����zءF����~I�����a�R�GtjX}����=����»��&$B���=n�� ��6�) ���NY���`���0�.~m���͟��y+ڽ���/ȹp�����n	ԥ�PʪL���;\�����L�pU�\LE#�-'��Oʯ���JKJ]�_V�؊K+mpx�:��ml\q�=A���[����3v��ΚZ[����N����Nol��d�^��9Y�V��VRX`)j��#�`g�0��f泊?^ IjB��"�Y8���y�_lb�C��?����뚑�. +# L�s��D@8͊�KR/�"��w*L�:M��"��\}@=4n���4c�p�`��K��A��2��I�p$T��䘍��盱��l��̴q��ٕ[�XՒ*���V����j��նr�
Q;��e��,3+�����=� �/J�<R.^�Q����J�# 	~T��p���n�38���x��(�%/j��[琽����>#T����*�-4���P�6�� �~%�ѻ����;:P�"���������?n�_�> K�eQu�\�	zF��r��B�o����7���Vq/|�8B1EV�:���|�U���'N��%,�n�n�OVv���I����,q��-7/W�y��]RR��2j�Ϝ���F��v�������{�䉓^�9
��T��1��##����

���EK]�ݞ�tI��FӦM\H�����t3o�	O���q1� ,z.�( �sn@W�Օ���A�z�������pठ Ӱ��׹8Z�zx���\+įR���<��ͤc��)\淑��a����Bw�����t+.�W��Z}}�����ڵk-_W�/�����DCy���f���,/^ly9�6""�Y
��@��Q �3;�Xx��nx׽�cNl�~��<g�l@?�T�Ju���z�B��.i��[Ir��ý�L^	r��w��$ 7� p>Hó��{h,JR~s ���軹o�l̇=�]l�=�L���B�
�8�9��{����@����砆�������
p�yI������b�}x���ߐw�y����q��a�*;������c�b>�X��6}�SI&ZyY�3�+�l������"o��Y�
077�Vɽ���X�;00��%8CîcԷ�]��
[ ,Aԙ%�{��8M� �����o<Ε(�^���Ԅ�����+��ޒ.~<]���� ���y)�̌tK����\������Yi�+1#+C���\��彂���إ)Ձ��e%K>MOcw1� ���ذ�4���N�)'A8�2R,/;ղ�2�����$���.��tІ8��l ��U��ܕ�*P�rs�-G@��x
)Qs ���I^ 0j"�����}��+��u7u@3L�V�p����9N�zGϤ�X��������/
W� ����d�:q��B����Xݒ&�E�����n�޿	W9]�>H/��Ï��-�saa渽�e�����
v�} &܈+\C,�V���0<����5�7J��5����~"�X��ٔw�Wvv�s���TƊ%�Oe����q����k\r�����آ�Jۼi�mټY�H��e���/-.q�&���R�i��d+//�y�,8a:����p��Abb�d'�~dl\~$1{��d�>O��ӏ�q U�\#���T��I�)�؅���>݁݌�23Ĳ�S,3=I��,����-=E"�@��BS&�N^N��e[~�z7�繰0G��%���_n.��*pe3q�S�Y�7
��J�����j�*���z:�B�8ǩ+C���9�b��2E�I�J��}<�)k�F zB�P����Ϲ�Y�' �Z����&"gs
���[=�  �N[܆[V��d@=oa\�UD� G�� �.J�'J���l�} (������w�����?|��_�o^��/���s��l�B����}�^�.�������,����.4��v�s�%��;���n��ib��w��H�D��
}��Z{G��)_*����W�Y%�c��d[k���*��}�I[K�՞;g-MM���n�%���&�h�"+*.�TF�W�K�&�UҬ�D'��36�,��$K�2{�+�sa~~��#������ڑcǭ��W ��D�iO[��w���`���[o{���7��w=m����r^�F�n���N���V�k�s��!������eC�6�����������A�Dw��pБ&��eN[aN��dZVv�56֩Gͷk��֊����$P�멢�wq}]`x����	`�b3�^�%�ع�Fkli���\cR>�}�F�J�Y��:ޘ��OH��P���x��P���0�DQ�D�����~�x�,"���;��m� 	�����=	��J��{O
�4�%}si���t���n�=&r���7��Dn��c�7z睁��!^F���r����y>�{Y�߇W��y� �-����� 3C�� �q��qD.�s�A�x�w��o"�wt�c���������	���MVYɔ�Q����cǎJ��_�����S�����ۍ����G�U`�
��Ka~~�3%�%V&�����C���/[Kk�-_��z���$����F+�t��7��+?1z�����l|��oBIp�d�k8�LƓ&�lb��R��-mf���Zl���&tM����q�L�u�
3���S�4W"����o���&���V��X���TY�ўF�s?S��^���`���C��<=$;h����ᴝ:���(-Jd���f��+��T� t�UUU>��A��**���<�`0쀞��e��6 
����!"҄�K����� ~� �4&����X�Sk�sV�g�>#���p� �s�
.7�d GA�3�Gʜ���������{�O�o�6�l\J^R
��1� ��:~u�cdy�tΕ�l����=��aQ+����Vn>/|�=���ʔZwP�[ ϐ���Dy�;��-���j�G�u�e4?�O�u���m��Ö!�K�`kHժ譹�ў�Y{䑇m�/ؠ���˗I,3�`�ِ'�3�g��9/�}y�\��;=.f�A���١omt|�G��v�q�Ϧ)�
�Z�0Ç�*�$W�L|w�O?F��Q�P�&-Ŏ���o=�f�[iy������b*(vyO����-� K���%�>Hǘ�����g�}�>h�24��E��� z)�������������F�W*��:���n;p�u�YNa����M��%��~y�ĔU�>ۺu��|��������d��׫׎����>�A��!��۱Sgm*!͞|q�}�[�Zvq��UZJF�N���������q�\�����@�FEy��]� �8d>	L�yV�a~/�#���G6<8�9��㛒�j����N*5s3U���@���z�c�����Y0���"�~�C����/��Y�$~'w�������o��g#l!�s����P��=���`<�g6E�7�b|z���<
�8�7R�
S�q�8���ѕo��	yr@�Ã��������K���5��b�V�<�Rf&l��U�7fC}�v�����?��V���^x�I{��gE��.�o�|��|���P�`�y��V ��r�&�loX6�m�٪ի��[%��K:근�<+Q[dӢk7��D�����kkh���b-��E�������m\�����?ne�y"�iS���t/��b��� ~�� e�P�����������l��U62��G�P�V#f��= �0�<J�z��0(��y :?�ء��@0	�K�TfY��ƛ��(�g��/�m��S����:�&m��k�_���H�U&����V^�e�O����Ʈ�����sMh��Bb���������΂|
HG��'�Cz��1�?���e�YA�K�̷�q��
\�@���&U�p������3a�5��_��*��ۤ:���1�Q�:5�R�f�p����zz|��ё�����:���LQ�үh��'K�4s�f�,�N8i�j\��2���fzZ�7
�)EP��r@=���N�7ō� ����W�R�\��lHq8X���[? P�£���ml�������l�[6������n|���	�Cؘ�H8�(Í:A���_�឴?��ҹ)L�F4��ɔ��6�ߦ��h;n�����Zvz�=��#���fK�-�*��뷫�]e+�����zkknvnrdhDt')S`�����]]68�gc�>Wuqu���ٰ����|��c��2��+���-����e��4e��|ƶnXm���>�t$�!3���Q��?���nL��Ȑd�CgRXX��0��N(q�W�!J�>BǨz��l?��G��jlP1��>Z���v�1��sV|��D��-��9�V��b�������2��(�n�z�mZ����QU>�0�|��S˶��Å+�������W���R�jR΁hcc#>w���C��}�1
Bb���Xhl (N�GcVy��a���7WQ�X�2Ӎ�FG�xf��zT~�GD�"�	�+u�_N`�P�n���r%-w�p_�M�t��h�@�K��&�C���c�ٱ�`���dg���3z����y7�gb@6�*΄�A��SC�8,�S�kz�7|��:CXc���&š�+M��";����{wj���?�n�$��YI^3cs6qj$��};$��_��@&I���F,��߫,u��ӣ��ϯ�OM`k�	Y��q�Z����}���[҃u?�MPN���NXi
3=QLO��:>�o�cC�V9�SQ��sMW[�e��F��8n55g|,���P�4-�D��@��]����*0U��'�Ψ]��J��v�T�=y���v;V�����RS�����H��GE�c6,��W�́f|�ᙹ��?�\��R�����gkm�k�zqqh�j��*��Qu8(���y�~%(����\ =$>#sq������4��IML0olܹ*�?O�������g�9�����:��4���-+-?k֚�O٭��fWm��228�1�=��W5����}?&���}���Lr�=�k����li�%VX��ҳE��)���]G_�
)}sD���8"�����8�ӣ�0��S<��ca�+'9<8 1.ߚ���ǁ>��H�'>@a���Ae?==�%���պ����e��X��F�����
ĕ&DbT(�se�K��`x����~n��!���Wz�Ez����1���BQ��-̈��v�.��Hz)^Ω"�E^�BwΞ����;ry!}He!��	�H'R��H��W3L��vO����x���=��Ɂ2aM���IuJ�YI��7�n���$b'۷��U�oht.3���&�ƞ�.KU��**,G������(;�O$t�II�Ν���7�b;n��Z{�_��}�[��3ͳ�EKlR"��Ѐ&��Xg����[���W}�͢��h<#��J>�����`b���5�H��9i{��[��5W,�m�U\�,�R�|b�4P�j_nM�Z�.�^�����t!�}]a�`h���G}_D8#�
�)rr�}��/�G?�n��VXT`��V�;c�lYn����Rc�ܲ����̜����Y������o
�	642n��u�O��۾��cV����J[rZ��HC�,MG�OLJqu ����XA�$r_� �#�N�`���������9�}ݪ�)���l�2{�[����������ވ�U��I��&�����u���M�Ŋ��dn"���f���DAR�p߈�/͈P��w��`�fa��]�6&r���
r��ɉ���0�q]�(Sm�6���c 8�3.C&�O(��Ĕ�ʁ��D�%NS�� �JO��Y�w�N���^�F����p%�x^V� bU >�bul�
7~LZZ��9@�;v�e3ٝI^��uw6��Wo�_������
�ʗ�`�N����KU'�IR�M�,n�E~R)��ѱqtu]J*��9�yB`:d�%v�u7ZRZ�8zƾ�����k9��6�|"���dX�DLv�ڲi�mZ��;�`= )Ù�L�O��̿:��	y��|?&R M�ç��;O<g���VU��2U�^*h9�DnFgC��ҕ� #|ND�ġa�T�/qQ?΂a�~c�	2H1"��OC��n[6��%��ĭ+2q:�YJ�a��~�m��k����:;-7sܶm����!�m��뮻�n��&��- {n�׋/�?X�ab H;{��бS��?l�>��^xy��.]%+Wϒi�c4v8���q��e}8W)PP#�;p����ɤ� ��X��f"�tq�,P�lW����n�f?���H5a���g���#����Ԥef��-��M5�wm�.*+�7���}��@6-�	��.�@���j0�K �^I����0^B�B�x��?:кX���n���!n�%8b�������(
����\k�9ʌ�H� c%`���322CG�+N�_e�螎%�m8�1Y���7���0�xFF%�G��ɇ�Ō%(�j�����j �
�t �AB�R�'YZV����}����ŏئuWؗ��;|����A+����m���2U��Y�VTZfee�*�ikim���~�m��fɌrh���̜|�IL���Y;t��54wYNA���=c;v�d�z��|p)O�e�6kΞ���^��-;�e���B0�/����6q'�t�*e�i�P��8�T]����bu-]��4��PCv�G,�,�Y���W��E
s\D��4zLD2B%CPq�b�i6hI���UU���z��{�-��Qmb6Şx�������Z����ww7[jB��[Uby�S6��h��o����JKX^	�!��b��Pi����Hhh�8��[��IU{�}[���&+�Xj9E��ő�(� tW*[YaT褔F�i���U*�č�h}�=�G`74ԯr�t��'8��F|��)PG����)1����2$�d%K�o���s����>��?aK�S��N�=�xY������ ��Y1E�%�E&*�W+Y�_h����BP#@K�A�8��0T&z7��y��s��Gy��5� �t�_����WR�o:\#w�L�^@	�#�������q��/\x¢c
w��)Y:��C�-�9+'��8��f���'�y��^��y�!;(i);7W�d��UF��Yu ��d�\��I�p���}6,)e��0"K����a��9��?��im]C��7b#�	�;��j���I����U߇tfb���;_xN|�����)�wH�<����@J5�	�6��t��}�v���R2llrֆ����`�dPV���̄�`r��O5r�Tш�|����|��bPX�8�^.�͆���?�k�ޟx�+��Yg�R�ѧ�����'%��d�����"�Ѫ+�lyE�	X��+�-oy�-]*nZ�O������,�;Ww�N�������G����Q�*����E��ž L�B�T����U>��Ի��3�ydd�W� �B4PL�!tr�_U�'�!ګ�Ѕ��$�������n��}�4�Hd��PG,+?_�:2�^���F�Z���/���[7)m3�Pw�J�r��g�xG�Y��V,�����X��� ���/� ���9�μ���{�K6��s�g����3�!K���8�����>p�a2��6��*�@�2���0�����0����=�
��$�}����~b&\��:�2P|���i*˹�����*���i�ю0�
�d@��,D�{ṧT�}�F�Z�꺾��::{�-A�b����	���&�]��NˬFBj
G2��358��xD��8��3bS�i�.>�.-=��\���z��>�<<�ccÃv��	����z��H���z
�ȿ��#��03Cm���hq����W�5�?~�+60�he��m69]fԁ���=9�L�9e@t+�#K�^9�W:D��8��/�E�r�R���;v`��������[}�*��R�쑧�����o��m7Y��j��04��K�+�m��������7���#�!��� @���������9����&�JWL `#�Mл	P� {����z;U�h����X@T���<+(�����ld�_�7�HO���SMK˖t0��&�!�U�_$1L��!��;!�S��ϊpggR�ю�����@1�
�3��b*U��MQYR�)jh� �_�i�#
iR�|�5ם���v����K�z�Jknl��sr���XyG��w1b]��������:��w�8.h�i��K�`l�PO<�/����m!a�H,s@���	�
3=�͛=2��Ƞ�X��H��Ei`�����1��E�P��&�i�	y���	��l�g�����YDhnA�Q���.���<Ѧ�f��D,Va�]e��M�E��&%�UX��T6ztQ^���TD^� 0�L�#_�_��$��IHU=(]���K�����)�@͑�Hе�V�Ǡ0��of�4�jG�U�|�^���BUVQ�Ȫ��:�=_��0��q�- ���Ti?p�����_���d+]��F&P���L��ﵔIz(�=�QI2=����Ǉ�!b�@v�JI�R���.���X��j�y�61�f��ʿ�?��ٛ�ل����S/�����oJ���*/S<TΘMM���
w�K�<eWm�l;n��u|d�F�¼W@B�ҠK/
�u�H�.������HGu:0q���yJJh'�5��3�v�\�Ҽ�ڻ���|��K6�ȵ嵡�Mw[UY�U��v+�L;z쬸�q۴e�U,��ֶN�g����z�)q�IS���&ζ����mb2Ke�+��q�f�n� �"-��= �n��O؉+%y�J�s���>_q��O��]�}��H<DV��f��엝�d��0=&�G@*��|�ga��8м������zﱿ����ROkl�c ���{��[���`ui��1D��4��}��X�4g��gi�C0�6�4�*:����zd�;�i�S6�oP���(,c��@f�ÿ���1���x��%�y�fߩ��2�q�x�/�����~���|���6 �^������ճL�!O�)�}6>$�H�p�+0��m��=62��5qL���ۚ�w���9��qs�)T�0\��h��>�_���f�2��)�O�v����9+��2�}ȳ���f'��8W�m�u�C*�˳Ғ�X��H�sȲ�����2CӒ�Be�؇���Ĝgj��vB\i}c��7U�ͱ¢R�H�hn�B��?�η�;��F���v��ت�����n��*���cw�u�]}�v+�˵}{���@�m�r���Mw؛�|�UV-�ں����%��RY)}�H=ݤQ�G�(��OU�qm�#�� ��Rz�k�꼻�f'�����՛�R�Po������}�߶���JL�h�Qd�q(@]��/eC}\�~/��|�<nHnH���W\�����������们��U�c�0�\|�7?/���]"��~��U������w��]]*�;�_�q�p��C�!�tZ�n�w���-'q���T�^sr%Q��ꆶ�"��)��k��|s?��΃	ޓĕpN<S���TY΁X����d�E���̪ˋl��Ev���qu��X\j�bK徬�Ė�_yQ�e�����j��ؕd[IA�eH~ ���' �w�
k�]��AH��Y���x�MA|�R�<Ȟ�~�c�\��ٹ�u�����3CW�>j�N�68s���觰���k��pax����5��Y]C�՝o���q͓���-PKV>8�q�Z��}۲[w�d�6UYqq���ں�k�~ݺ�VUUn��zi��\��V���������7��{���֫l��5���9��2�Pf�X��M�P��+D@TY���Ib�*�]��i�|���m梞W���OK7��d��o����,�j�s����Pg��M��5�����J���;�KX?T�eY+����ܿÚ�HIw��b�[p��Et�n#���U�������3*|��T_�B���ka�P�L�}]]������ Y�����*�bĲl��~���0����7h{��w�r�Fۺy�m�t�m�b�mݰF���VWW�浫lÚU�rI��[Um�7�����&�W��+�o�*[��Ҫ��r}��z�D�bK��3��SV?����f&����{�[�r�遹�*;S�nO=��
K*]%0&����Qqkbw}c�����Wdsg�
��(�����)Ѝ�F��Ā�ϝ҃N�� Ϋ�n���#�ő�Z�D��nKLͲ��
�g F��yw{�����_mEy)���8Վ.{��GlGJ�7.�&�G���i7�|�mܴXD��Nߐ�?p�:;��t���c�r $���H�Q�˻y�c
VE�r���������o���Bc"��%K:�S��Ԣ����}�]�zE�O�aN!�%`z)����#�����>���!����qz��f����0����������Ս�����q@�^�{������-�qu���!�<ٔq(�P���k���6|���JWO
L{{{��:|Õ��6koow��߇+�Yx���wN
�d�.C���Eى��L��ڰ%ΌYEq��s���2�m��û���h������Qw�z�jl���Fe���Y��#�|�w6[Nʌ�\\"�]fk�-��p��ٖ��F��s�c�Ǎ�EQBs�E2���D�8���F�U ��r�:�Y֧3h�$���x�ZZF��r���s��u!�peh\8c\ �  D�� ��8���E���9 H��
 �\����l��V#��K '���إf0J�Q���������޽{lDLy呜h��v��I��?'pb����^۽�;|��Q��}	��H+;��
��T���7"�8���w!W�*X�����;�=c��2�?g���nq���D��P޺�領Y�<lڴі-_�ЗG'�_�.��W5�~��b���`渤�x��f.��k!3h���Um�/m)H�a'{�����y��IV�gdc�tV���P%�8tUؤ��-����Z��~�ņw���#�,2�n�2u�lk�6]���p@`�m\[���ŏ`9r�9z�jj�����ϜYh�.2��R6u�4��j��/?k;�~���oM5'�Ⱦ��������=����w��E{mϋO�K�>i�<�m{������?e{_z^~����N�8jC�����Ox0���Ѱ)1�y��̫ �%���a�-8P6��k�I���+���k��s��;<)��ݞ۹�N�;/N��� hX/��t%���#wY�#��U�
jpx�^9p�v�9`���[s{���	Բ$��)F��H)\`iy���4�+{���0��*w�}dx�zz������1�=]��v��;���|f#p:��'E	A'l�.�ޏu���
�_�3�)>i�Ъ�}��ʛ�O���n�-eM~С�)�OU�h�op����os����@v���N����?�Ӵ���o����B�ﲎ�
ɯ�(���zl�A����ǀ�&xsw�����n�-?��ӆH� ��s*(TjHc�P̴.o?�-���Du��S�l��}v��A14�!��&dH(�h�
Y�,�-Y�^Nz�U��ۖ�l��m��ݗJ�_k�^�ɮ��J�q���7�i�z�>����ضM덝�O>h�=����k�9�Ϛ�}�����Q���{Ɣ*�Jy�{��Qg2�Ax��)�4p *���
+W�xb�:UgGΜ�ޑikjﳝ���3�6<:)�+Z9&rϽ���i��Q:�Y�0uFi���;0j{���{��ַXW���N��Ĭ�e�Yjf�Ү�đ*�0^ D���%�fB�Q�-��?� �zz��{��gl��]Yq�zf�!�B23TFp��x�ƺR�~�`��G�C��P"_��`�1��i��s��1x2p�L��������7?Z@���l�*�U�zw?����";w��J�k��խ�]�z��J'M�̸�mԬܒH-����~u߼~C]��ܸĤ�;E\�D��sY� ��MVv����Z�bCs���6�*�K��Xe�����0v}*��QC����.y���kW٭o�a��y��p���ኵ�j�rۼq��t�uvێ[����l���dq�o���YY�j�lRB�U"����1R3�S��@�9`թ0o  �WU�%Bg�Y� �G��f�d�e�ٺ&ۻ���8uκ��%ʒc�q�{) �X���� Bp���E0&����v�Ǟz��:���HlF��4q�I���$���	xXҔ�<�)/P�¥Rt)I���;�c���8����׷=c��I���RD,k����F�V���������q����+`�ׇ�����fF����B>,�d��Frq���X�^Һ��6��dl�M�w8w��Ư�s��B�ν[p�]����,ɇ��B�ܓ>�'�F�𜿧��: ��{�#s��s�0Ei��ցrP��"��nq���A���mJ~�<-�q��Q�a�8�״���z,%F9�.I1�O�6�	m�f\T��U�mh�e�r���p,�؄\�i���W&��}TZ��"�������`����ˊ�+,�0�F���CG��o8o�55�svWg����۷��ݶ�v��n��f��ML�Pĥ%����IJ4�h�Q��**2+3�
�Y��+0�V�f�M*y&��9<9m}�8*��m�ZBz���ipp�),�s�������˻�Ycc���	���|�,��@A?84\�ݪ��w���<v�z�1{�Yy����a�ǤD�l+�\f��>וUdqHb|6�R^i<N,D2c��i6>�Oj#с[��MM�ci����ã^H�o�!����}�H�!^�"��Q� ��Cj��F&K��dCΝ�S%e��_)����)\'Z@VybR�����k1��%����!8D7�& &R�b�D�3��a&j��F��f��(.���Z�����9oʐp��1��������.�_`�В��o��3��:OgC	��ǜm��:<��AS��Qe�^��뚖*�B�0B2A0|W��t����X	��2R8q[���S��KK� �4��s�r$����e����R��	���,A3.	�c�ݳ���6*F�F�3��3�1c��.4�%��2.��B�B�T��|��G\B$��k��9�i�8��6Y��yL��;�/�v�FԘ������K��JJJ}�&ӕ �yZ����oC�UᬌP��`�s�R���Ho�?ND,I��MR���}Tfn� ���FFm����>��|C�}�[�ؿ|�������߆|C�c�C�Va�!(��E`���W%���l����O��O?oO��:qV�h�5�w���vq��D\���, OJ˴T]M�922f�ij�j�gԟ�Jp㱉����, Fe�aݣ߆��|�B����T=�ѣ'u�w %~�>����P�s֝�aR��������,o�����V=@�_R>�c0�\��� r�/�X��$m�����C��l���l#8j2Ψ���� ,��u�Q�rNQW�xt�n���Q��)�z6}�:�,��~0q9ǆ�|��)/�!�g$"�P}�@�g���{�����v��)����9��Gm����-�8���[͹Zknn���A��Z]m�5�o���f��!���CL���I?L�U;�{�a�!1,_湻�Ǻ���]�u�;6��#�����2���߮]��}��%/k/��T��J��^��0>�	��տ��;~�7B�g���P�v١�������.�Uo���,l@e��N��x)0��A_FOPZVn�[}C�5�vؔz���kn����}C@*��4��Akk����&[�l��`�jz�'���%�`�D0��4�=��cQ����R��ٮke��>�F{���ܹ;u��&}#脃��!�9N�r���;`�[� ��g��CGO�ɳ�V��n��}��7d�|#��h��5
�=�o��f�N�I�U��:ScC��TgWo�dۯ�`9Y��|e�a��e�v�5W[Qq�ut�����]?�}�6[��
e?�Z;zm߁#��ڣ�m���d��e޻{�hi�Q�P�*L�q��K���#��ۛ|C���z���S%y��#�>���ʰ�[6[iq�Q���A���M��� X��A�L�^��C�Wl�usK�mܰQ�~���'h�� J�^l��p �r0�x(K���:���q���l�<��]`�#͔%�$�#$�\�	�ޟz�){��'����ZZZP]> B��#�I��z\�������S����cv��	�i;{��ժ=��r��Y;q�;���v�h^��Ƿ�`Ϝ9�0�����V�sg�9hs��ѣGlph��������o�Ź���ي�C���9����ջ��N�z��i��	t ��_�`���Ժ(ˁX�U���Y��zV�lܸ^�V#?�7

�,�E�D�� �hEF/��O�UUGZ<rܺ��,;��$
d�:�ff�8qfK���Qkm�����n[�|)�H�7��C?n%�U���I���z��i�l��8m�y�~j��Ĩo)'*�뜲sQo8���&��mjk��5��lm��v�t��?x�v���:��g�^=��=`m��=�6<>c��9��_j���N��Y��)_��/Ч\&�P9�@Mugm�ev�5[%���(�O>񜸌�V�|_}��VP�k�����3/�8�N�o�j7�W�')ݭ��/�����d�e�ۨ��3P��nJ0����� �ScI@��o{�=V, ��S�(���m���f�'����O@`�pH�:_x*��0B*c�=��ĭ������I�-jԈ�ppp�!鄅	A�<B���P�{om�}Pm��¤S�Խ�é��/��ǏT2.:7���A�Xii�:�v����P��L�a"9+�jkkX��S_[�η֚��9v�C�s������2�A��1����g�tw�#en��hkk�)A���2��[���m������D�j?��}�'�?~L��-Q�_�v����v�w�V1Yb� x:�P*���^x{��R~/ �
~�KG�)�&]=5��~��ǜ�<��>�����%��a9q�
P��+sD�lK��]]N�DN��� νf/N7D�dc�t��
 ��DE���0��;,e7*��|8ҙ)��������x���~�	{���f�?�ۿg��ל�s�A�v��i�Q�|V��Y]ԃ׊c>~��N�QOz����;n���o;w�C�j�C�5�I,���!5��lK�)���Ŗ]P��GN�m�R�3]W5&.=��ݥ˝�V?j��!PZ�v�-��Ú���=�z��\�X�'�!g3�1KM��E��j(�Q�UsU]����J1�Gd�p���"kqI���O<!N��.Υgf�C�tо��t½�G�/� P��H4]�z�-Y��7�X�|�[6�@�F'�͘�CYBϱ{ K��E�d�Q2���mQ��᪎��D��1p�֍.�=:i5,�˪�}�f�}���V�:(�.�(�JYHT-^d��VR\(����
-?_��S�C�ǝ���{�$H�u=ge�(|u�iH�L���̌������Iy��
�Xe�Ta[qq���XQQ�-_�D4�R�j��j�2#�����l����M�9Ҩ�uJ�=v��M�W^�r�*���4�R�T�F�H>K�R����DDl��� �%�Kr��޴�HO~k�7Z�yq;��;4bC>7T� Y��( �;s����b�
��NO>X��2`_��7,G-:P�=�?2��]�9g���Q������f�n�b7��[�b���;��4�1{�z��|���Cv��Yq�mzn������خ���][GmtL�߸@2!U ��<�-��#�Qke�yPiPɌ�'�/����V�Ӗ!n���&��믲�bu�gV�q�
�~�6[��J�{�}�	۳�+-)����>�u��V(�3�(�uEF���OY��o}� �cQQэ��5<#K�OO���f�L����w�8�<�H�v[GW�=#�K�#388�������6���.�Q��i��]( �H;Y��dI�-[��uwCCC��*��Yt��7��O��߰<���)t����,N�y�ǖw�:�P���tq�����5;zX@�zs*i�M8G��ѡw#�R[�!�wNsH�kOw�wʍ-����zu,�M�����a*"��!����a����o8�u��e����^}7$)O���3��=��D~�a�0�K��ɓ''%�s�y��e3Q��D{H �����&Qv�����mQy�uH�=_S#M����rҦP��#�f��b���
������+T��V��dgjꬴr�D���7L�	����NgO��n��6^�ʁTAy��~S Z$��@���F3�S�R���I�@����l?����o��n�q�]��J�����r����uk�}����ƻ}�\��T���������(��N�/���"�{g�YQ�b�-(���bK��W�e��Nupe@���|J�ڃΰ�^�:����'-%i�r���+����FHiY��Z���*��?�j�%J�Z$��~�]��w>�޾\�QH����/^���U���#v^u7k��y����i\���P��]0l�'��" �S���~�k�p����o��׹�4';�uy��\��(Èǀ"�W:iY��}�		Q�E�%KŝV8���
-$`�d '�3a.4LԎ݂:�Z�[G��q~�8^t�0 p����tD�>\S�(;+�XF� �n���.�#b#����������c�$�e�U��m�:�7ܶ������>���n�ֶn� ��s���R~�L�C��g���J?Si�"ي2�(/��Zy�n��A����U\R��L����l͚�V��}��T7o��z������`~��4��9 ��������ç>-Q-�>��ڕ��ىC���g�r����"Ved��q� �)Dv�t 2�]�Q1���3_��}�	���Z�Д�M��l��c�jA�8܉~{�k�j����zǛ}�>�<�Ľr�����ڢe�m�����H���>;up�=������|P"�8,2Y���5�2K4+ZCS�:tЉ!=����;)�jr�W�!��ǜ���V��*4��I���?SH�D�""D7�x�q��ϮWl�?-N!7+�ʋ����G{˛���K�KJ�+�����3������e}݃����{���Z!/S����c��_y¾���mb&���V�N��'�x�X�#��d�+gؙ#{�HE���[��\�U������v���i?����_���se���� l��x�B-��2���w=�$#����j�/����S��֌x�����]{��9�4���q��EG��Iw�Nޠ'�וb=⍹LJ;ހ�o�V��x�kl���\�0#[uI��++	��$���X���t�� �.YB`ޑ�G{��C,V']f	�;���e�X��X��y��$��)�]���=+z
��t���ǖ�-^lݝ]�O��O����7���ʳw���v�ͷ��?�q{�O�����ڨ0���#��;��!��lT�~T�����R\u���z	���^�8��Vq}�N���`��o�����}�^���֮��M/,�H7ʴ 
 LE��P���* _vPb��c���G��|� *[��~��Eߦ� ��M�[c�?��#x�UW��U���$��!���Q������$Z�(�i���Cvݦ����|�-[*q[�P�hm�c6�~*E�C��MOJ�
O�kR�ȵ[U0ꕓ����={���۪W����"�*(��ب��#&�̖d��5�*
���[y�C=mi�3R�mF��������S�`Ѐ�Ll�����4؞�'��.8����ڑ����o=m_����T����5�rζ��tu ]V[�h'�4ٱSM���S�NH���̬Bџ*_���$���t5bK��Ishء�'��e���s��16̖�v���#��/;;�8j���W����c[7_a�#}j�]��o�WĀp�S˘w	w��2�w������&	+7'W��:�Q���=/�!õ��#� �Z���S�]0�bN-\!�p�XV�qⶋ��3�?`�����2��Oa������e	���["y�uʺ����e�t'�Kfn�b5����a�-��-۶�*q~e��JJ��P���#�@�='��1�����)H�`����\��&f(5}�8_�M�MU<�ٖ��_�#��	��_��2ő��Nj��6��L�~��������b�֮��V�Z�Nl�O�ۡ��l�b���`�+�����<FI�akN:�0�:c�T9µ�i�`cg���W��g?�E��d��w�öo]a��[�_��/mbl���-Ϊ�hTV����]�����~P�'�cd��w`�=c'�6X�����I�o�ː�8ŅJ��7�����q;������]�}�}tOe�<q�>��߲�W\ey�*{�{�����G;���߶_����{?�!˗Hs���>����K���M������ۭ��ع���'����'5�����*����3���O�f~冭��]���hMN.��c):(��Y�`�xLp2]�Ġ;�� ��
�S-���\��r��.�G?[������x2Tn4�Q�RU�rۺ�j����s5���&pd�9�M��*�d�v:�RK���s���d�) ¾�"o�VW�E���͙ީ�a�[��VKT?w����?}�o���+%������ҋ/�+~���o�~�'ޡ��lgN���2}c�$$��������Y��L�����Ç]���촕+W�:��m 2L3R��< M����:�������� Ʈ��;ub���7_Q�u��8]���a��D��l�\��#ꈙep���{��>KQ�a�h�7�D����7��y�7lG`��FE�O��H����2q�A8m�`���F��Y�q��z)Ke�-Sǘ��Ïڧ?���u��\
������?��OZss�����U鎊/�'��h�F.�Q t�Qh�|�:�+���#�@�G(۽������@��~Юںֆ�k~�˟�ڳ'l����aV{�B^�T�0� !A�l��
��1ki�7yFX�!.���9c����R��)���4[��Һ[����/�g��Om�8��D�B�@eO>w����߰EK�,Kl|rTb:Ǔ�ف&����U�펻�I�s�~������ݳ�V\��6_y��Tt�U[�m[���������
�r����e�ރ]�����T]�-Y���rōJ�ALdEL�8i�YA�a4U��F�y�IOO�א)"
���3��t0S���Z�@�d۹,�S�du�\��hF�팋#JSYT,*�y��{;�$1�ZGK��
L)���	���"�dq	��Aʴ��+�{v��zaV��`����7oPcJW�F���V`>l���?؍�o�� �3��DD7د���ۃ�'��ץ&WClX �A��g��QØ:#ՉʈΣ���Ey�Y�\���*?!�a������eaQ�݄���e�:�X�� ��s]��`�b���d��4'0��6aP<Ja��qC��%��d�z���%U�e�V��!��k׸ȉ�^ZZ�u	'��5����ԧ-^\):��ƆFklj�9�p��I(}q���?V����y}������ 6>M�9n�8e	����|Į�~�����_��_�S��|Tf���B��UL�.��,Fi�~�4�c���U���ы�m-v����߰ΧQ0R������������άM�f��a2Y����ڹ�����MYN~��3��̖��plo�@e|h�z:Z���(B�W�&�3�� �;��'_���9��8ǭ��ƖTJ�[�"�ٳ��_�e6o��bś���С>�nJ`��SO���;��U�Ȧ����{־񭇭���J+�H|1��{Ȳ��2o@���΂�ig�}L�[eA '��-�� Vp��N)�q>%E��(?6��X7U.vp�x���H��j��
r|�KAA�/����QG�:�tub���q/gk�N���a��u<#��^"��'Ǉ]o���>:�#*`�x�6o�X�z��wblR�g�}�_��粲�'J�~.#��r�_V�.;,� `0pG�c�E���ܹsv��i��)�_�c�G@��,\>��k��Z���G�)G�zi&��-�K�-(`�P�[t��_ii����.���lQH�"}螗.]�~	�MojjjܝN�lV[B5��������Î�8a�w���|��������bBސ�&��D������bƎ8_,�<+�����bT!F��	����W-Q>����˼]F�o��F������m�@�j���Й�t�a��7�́Ŋ����������с���z����#�,�hL BgeJ�K��W��Q;Te�����%b��GE������
����b}*�<�] ���ez:ڬE��6@qQ��F��
�u��Şzz�-^��
����'�F����
�S�Mw�fe�ޠ_�H���z�%N��$�qv�ϫf���z��޹�3�]�կ=b���l��I�T��B+q
p 36"���#�O�3� @��',C ���# F��6-����}=<�)QnIj�p��FG8��qno@\3���!EqN	����O�0�Y�7�� ����N��n�Tj��S�h&-ivB�)�H���h���Fy����*ݧ*ܲ�|���V[sڎ=d�v�l/�|A��i�m�[�r�S��3��O0W�r�\��T<Q��򴵷��J�=5��ce+p��x�U(tp1�HNb����,�`�)���A�	B�AI'�q��7��tx��?���e�1I^��t���.� �::�[��ѕ����7S��+f$K�(����:/_Tx[ZmkV�Q���D��l+,,�����Ze֌>�>J�K|@�6�MU����ʭ�/^��Ř1���E
�1����43���^�H��2!��mΩ�(��-@*i�ͤs�jF�s����,�M�w���>�K���|�Kv��+~���׉%�EJ���-�σ��G��@+Ĩ6 =)��Z_9t�jϷZn�@�$��M	Ds�� �Ο=n���o~�m�-�:�:�Y{����~��ʫ� ���7en����4s���?!�g�﮽�����ٚ:[�r��UZ���}��I�q�>�ܙS����-{��#V�t��W��ش�+�i��ş	�R�wF����٣�G"��
��<9���7��� �'��"i���V�U�����Q��bWc�>b�8��A�����B�*�68u�O�����(�� �G��;T�w��8+D]���a0��R��ȳ��$���� �~x�Oa�M��K\	����G?�Sj�w` l2C��G��[�e3H���Qgpj$�)��o8�0��5�,0`38U� ��J�✗�$@�@��be��_ew��ix�pz�����b�"��r/i����CZ�)��I~�+�f�s�I�#A?0%�����T�-�]-��jc@��ʁBiwN\6C ��Gx<�.$�T��y�QD{�������v8�������f?��`���w{��e�����^W��q�N�ny&}��<\�4�n��ށ��+�������Wm69��%�m�֕&��v=��5֞������n�W�^�*z�.��`��	ZĚ��\�,?#db�v�;,��Ѳr��A����XQ^�՞:j'�l��ڿ��7_���7?���i�+)[��[�Yg�9l>a����b��q�D�D�������/}�k��7�>�<�=���]����{D�g���7��g��s[KW�u[^�
*%�F�@d"��9� Z.zMF`���*�+��(eq>m-�4�LJ���%0�
�Y�gFwY�UR��Z�$u�$��L�l��'���=���h���5XWK�������k��Yq��%0#���93jR��>3xB�!�� �#]Fz`�	�1��hȾ�^����UC�Vx�ֳT����rV��������_/�LܲiVV��c�9n6G�k��}�F����\��O=e�o�6�y�G��].��!8���6A|�ó;%\@%�������0` `L � Ns��.�.퀕�G�S��
 ��Kz�U�,�F��S�F���*̰g��]~���/t��6����ZYD����'~�XHP�����9-d&�>�� �O;��{���~��~�W�����}T�;Ĝ���سj�E�l$���qPV��L�㲿LFi�w ���)�SJ��ۧ��5���{l�V)�Ь���F�!�f�r�c�E����.�0��lS���^�����Po(���g_xَ�8�S0�%�[���L`�Xs�N�����W(0U��l�=s����������ew��A��Q�vٮǿb��6��_���˝+ݷ��}�o�7�d;n��::�$������e��=�;Ϗ����U۬���k�~�Nמ���bd�%q�웊5-�J����Έ�{z�J���}�6<�i����j�L������W-_���~�u�LЇH�1���ؤ�Sb_w��g�	L���ӇliE�ol���h�$�]s�u�������ꄑ�>q���
ę���|b6�Hh�pLS"�_Ņ~
Ѳ��Ж�X��1�SO�reh@�i���x|��i�Ҹ���n�j����]b� ����i�-��������F��p�8.�\d˪�{^1W,_aK$
��֬Y�`:<:��ĩ�c(6�	� HLG�r=��5p}p�&��(����)�75�O�0����-���fz�b�ĉ8xGX�#��9���'�&�Ŝ(z����p�4�p֮� �#cnѪ<�<(��=�#X�?��� ����&�����g?�a_�è=@�����O<��`S��n0���>c_}�)QA�{frwV�* �_bf�̤O+A��&�Lob����v��qQωKb;���Y���v����R�TU@�89��=���q�>��?�-[V;�B2p���ه������;ՐS��Zf֬e�O�ᗟ��NqK!x�Jw��C��'�� �;z�JfF�j��bc�zb��U/Z�8k���C�����x�����!�5�g�	�%j���TÙ���Ȉ��wښU����x��6ة�G�ƛo����+_��}����[���?�I;~����*WY~Q��&��Ɍr���DGl��ߒ�F���]v���3�}�m�t��;{�>l�V���o��0Hǩ�cC�HǕ��K�ץ7.��噑u����	��O)@�esm꓁@f��j?bjin�6�ĳj�*���O��'�Mmn��F5D�����./�pO����={��g������ӣ�`G���Z[Z%*w8hNH�@�x�D�B�\Q���t��G6)�S�W@+�9y&ԳD�ا��H#+���LR
a -1}����0�I��:+��8P�>�ep~���ꨰW a����3�ѩ�^�I�+4�>�0��=����>�3������&y���7����G��y^gϜ����J��&������`w�u��={�}��V��u�W�/�-|��7����D�I�����*Y��]@���/�%�?��ƾ���6��� �/uz��I_����K*@��>����4.�0�g�wv�Ab� V��X	D_��E,�\�y�G,[{S�Y��j�/���ۖ+�(�;%ob6���k�������e�����jep�Z[���P���R{�ת���8�U�S��F%�<���>by��W�m��*"Lq}.D��qDp�ܬ}�+߲W����	[ԳO91�K�j�s��U�=mm6����Xey�@��D�T{��[���G{ܮ�(Y��_��W|�1f.�H�fɬ�X��T�4���'dYEQ����ۛj���{������n�C}�CvB����l����)�I^/I���Z[���]*P�������
���Z��z?�D�����lٲ���}�h�D��CgΜ���~�]{�u�J�}�\뭷ݢ�UF e /@п�+�.�Q]�X/@��E����^�/�+�� �(�]�n�oǶ��w���t�Uh��J�r��H��xf/	T"p� ��%�F
��C\�F�w>]��$�+"=���0��f���[�@�{&^8J¤C���y�Y�#�΃|���"P�3��PD��$|ޱ������7�pw@'��"t¬���>�H���m�W���	(��ʕ˭�|�����󥡟��'�/��/���XKS�=��w|^��2��أ4(��M���m�n��.���@�8�����K��g̲
,Q�;�f�ҙ�qy�H#�t�D#�w*�4q��P�����"���"*F����?��Ez�H�&���ғ,?=�N9 ��o��v�� �V<&���ן�׶~�uV�l�55֊˪���%v��6���N@��p�Ϲ0^�����;T�[�\���Ƴ�#�®Z�w𨸑d�/����P��|x���!�z�,S�����S\Z�DA�cd�E��/�v�}�ʨʨJ��H('�2��~P��2�=[���&իw4u[i^�o������������,QsG�k�����O�l�pT��T(.�� �6zp&�D�8Sv:��_�5oLNg���X���]�|���Omٿ����b��|���c����C@z��x�>,n�jI�m�~��am8g7�P/�C`t$�{ʂ��]/�V~��S��pc��5k��ښZ�  *�O+�cr��!�R�����bm�d	����N�Ɔ��Qk 8�w�b�O<�ցZW�)w�#�P�#�h�)}�: �6�FEK������êt��uX�}�B�������UE�	��4�4���d�@�����!A[�e�	���<�������%��>[%��c��������s�}��}���`�;�7^^��jB�Q� ����wDק�6���%d
K�|w�)��D�z��Vv������'�����O��P	\�`~�2�$PT*�����c��f�b;w⨝9qȾ�o�d�]���o� 0�����ٟ���~U�����m�\m?���ن�+-A�0�LT4 n�iX�	��K�J<��<�:+D�|�}�{����*��-='�7U�Ы��MZ&F�(�z-Y������<5��F������k�#ݮ;,�KJ�|��9��Y �3���ęP�xM�����g�Ξ>e3/�W��?b[�ڬ�b`b��7��S�`�`aQ�8v��	zJ�4p�a�r�z������h	��2�r�w:w��]���

�����ŝ��7��u���K��K��vź�j��i������b�3o��HUp} ��={��|ȁTN��E�����ɓ����� ��.ګ�M,��BX�c���11 QިHB�5#0���*C�P�q�@Z��k���\����G�����>͛zf0�<�.����w@��.	CZI��qD�*	�r�C���A����D�D�T��0��g�@�䅓0hS�yN����꫷{�~�W~��������m���nO=����J0�)%�mlxy���	�GiPy���Z{��|����>;r�M'��'�*؄�LN�Te�g�
]�OJ��Ϊy�=�O�;ҋ�˳�]\8�^�Q2KHu��ϗ(N7]�����7�hki�7�}�-_��E,�S�H��9j/���V�Xm}�>��S�~�]�f�[2u������LSYpTU���bQ���f�d���b�\���;z�� .�l��E���Y�ɔ���~��!���g��H���u����l�{ϛ�0,W\!�w�뉖�����������YVR\`e�!Yl��^Q^h���n�Z�hkwT/�M�6Y� J���),�(.)�J=���"�[^i勪Ի��Y��b����DFF��]���d��Ï�.�C�cj�����ST,\"R�c}vV6�c�;7M#+--w�ޞ~{��|V~^d"��3���	�nTF � }d�O.?-�g���<5xcl��1�  ������ �4$���cP�9 H\�ƿ��b,��D�͹%�)���xp��=W��AZ��kDu�6ʔ�Kpr����Ԑ�|m��:Iv�0�����3�N��P��� ����m8��i@e'���7�r�6��Y��w�������O�cn)a��q���Ej�˨{�G�Moz�:޵�gQ�K�.i"�L&��Au�@��䪌�-�ګ���u���:��o?i�����_� +��b�,@��f����.�K�vJ=�Ls#�ġ��UF*�LE�"������"g�_bm��wp���������qp"T���=j�������g�λ�b�}�j��G��nm�%$���}k4�+6� D+++}� 	bb4=������9:�N�m�ϪA��8��2���	d6;e��66�g��T,���������/����Jq�Jupp��'3�}IMq�{Cp��9'č�r��S,E�}�ˏ�����sdI�����)+,�H/a.���<uJ)*kf�*_���=0���������sM �����Vlb�\��u�4��ڧ�cr6+���iM��l�Fg���n��Fşl_��l���%K��m��0/#G*C���Qɧ������o_�җ\*�Ymm�UW��i\������u�C��f�����U�%^��=u�!oH@�L��Q�Q!Š��{$%8Ÿ~�z`��$u�#�C��h��A:@��,5��� ��N?�b�� �v�&-�O���A�p���!}0+�Kn�h�4zU��1hZ�?�s?o+V���ھ���kjj���֊6;��t
���5�7���(����e:RJ�>5��T�s��>�Г�5�g�h����n_A���QD�\�i�W���Q�Btp�����N�
'���&�1�KE��+��x%t��ۦʟ����[w� �0�����~���7��/|[��[���κ��۟��Gm��6:4e�=�=��sN����q�Y���4t|��,������D<F�b)(S8�KrR�:v���v�yzr��'l\`��4�X8[����C�l�U�w�9���	.�	]	��Fe��^��%?��3���w-;O\�Dhv����G�e9�i��萸�IX���V���8�#N��F��@zЛQ.ppN�a
���cjr��/�i�
\�8ӭ��]���+����B������!���̒RH�❾�@*zT��P����E�"������656�*�k��Ύ9�M>��N���"� dq@���|�?���©vw�ګ�A,�"� Fx����������͉�Zļ_�$>��1���?\( �\Y ��O��������!��G8a��PNp��9�>��N��u�j�t �'�����U�K�_��=vܖ.��;�_u`��공kW{��������v�=w�`�c�?�Vq��Pޡ̃��~�&��A	����| �������O[Ww�D�A���j�����5�PW�ͨ��Re�S�J�RY�T�d��5����i֛O��sRū���~jd�&%:s��]���	�3ϱX"���+�mo�W"e���QXE3�h/��kg�ԉ�����Zq�v�D��;w�֞y�y'���\��+7[����j�d�i������km˕[|~����z�r[��R�v�-[Va�+���$�meE��[��*�r%ڏ�������m��b���2Q��*���H0
��h7K�TN�<e��G�5�ٳK��^�$V�Xn����/ﶄ�t�y�M(<6pf
Wff�ը��W�7-�ͧ329�%(�`JM����,%%]��&�`�Ur���`j��=��O�ALT���`\\YY����v�}o���S➳EJa*�HJ�2��j� ���ź@�����#ޙ0h����Y����ч����b���pd��Pء�g�pb�<��Qč�L<�i	�{,a����Pg���+֭�F�z���u�$�\T	�M�� PS��.�҉�8��� �H1����E܌�47YwO��'s�G�7���G-B< 
��_ye�s�ebP�r"��C.��/�h<�v߻�%���b^��2�]&b�Ҡ�~�އ������~����2r��P�wjF�*�ef36<�kc*�$5�L5>�,e5Lf:�m�� ��^W�#Н�*W g�B<L�Hr�Ζ�J
rm��u���t����Y����o{晗�^k/��]�y�����o���Ծ���"�6���#��ô't2+V���4 F��"q+lZ�ȣ��M�:c�3z�Px���C�؟�UD�������l#+��Ggu��}�ٽ����7�ZgFf�Ni�2'2~��_��۰a�O٤�_>�9���F^�9M����ҟ�.D�h�.�q�ҥ�؁��Ÿ�E�qQ��'\�+��"��NXIQ� (�u�4�;�]�������,��ɏۯ���ڝw�����m����U�êZ8�H��Ɉ^f�A ��|q�A�w^_��]�б��^��۳{��=w��@4��X�)'W� Z�rNN�so�K8{:"� b����8W1�#zJ��!�H�~�'�i|t�,1�~�8��ƌ8O�H<���W]%I'�9X�Ķ�����ۛ�S��g�*j�B1)�C�'� �>g����u��o�DQh�\L�d�}��? `�=���*AUDx�7����C?a�ٟ��}�_������y8|�/ׅf�cVJi#䌃���2b�NTi��g�\�e�-u����c���'��V�>%G�|��-�m�*[���V..���l[���e�v�b[Y��V,ջ�Ŷ��ܪ�.�����e��OvE���0,ٵ�����l��]�v�jq��z��6]�F�%��3s#C!��I2fX<��NkjnU�,��M��ڝ��"�P#o�U��n�RZ�D�v]\���]�y�o�M��3i��]��&������v^���K��&F{|�iz�ߒ��4�
��qw�y�z�B�s�)q�s� ���,GD�����뮰j��(/����o�o��`��� H�����x��V�����l�/9��3St<��&�ty��|�V�a'�)p���L�� �V�Qn,�7��*����
g����q��\�F�����=������	۰I�ZV��L�7�����m�+�_�l�8�p>%�A���e0�,���5��}���D�<y�ﮅ��%���vL��C�g��w\7DT,�\+��s�Ы�:�h����\�ðSk�a(��q�7a!0�{8�TI4ʑ6EA5��{ �l]�+Ё�FG���hL�b�z6Ҁֱ��s}��YQ�L��7��8a���KA�U�M�Y�ʧ�r��v��7��7��1�X�ܷ�;}�X�ѓF�ע6�s�*7:h��f%�9R h߾W����e~��	�x�xi�V��~h����IW���L�Յ�搚,���3����J//*�E��G�"��tKK̲�$�|��LKOP� ����Rݦ��^��j�)"�T�4����/3%^f�qr���W6]=ef�zLD'��o�J�(���h�\��\�Q�X��.�3c��&O-���9謡A�Y��Bű�9*���aV"Y���{��h�1}L��F���ވ�G�&�8�
���$�g��r�MK
7gܰ�ӱ�G�ܹ���ڮ�/+6�������0�������������S��[]y�H�q�|pceG7��Z���˳��|Y��Ȣ['�~:�Y�\�3;�� h��jܜ �����}��h��O����TC���%��Οo��(��8�'��cTʪ[���OaN��E��y�07��`�R6_�ܡe˖�����ȊsW�*��N����X�FeD`����F�w: Oa�O-4����b�'i#��">�����n�q#��L�6�& �'t��ݭ<�j$ ���y~=]�DX0�J�[o��������K�_���_��_������$r�O�g0i��6w��g� `�ʁt};�m�F@'tD�� �EȀ��}CI��2�B`���%�������ش�S΢K �q4I�i�a�3"q3�rgC�$��U��x�x�MO�p��9�rMԷ�Yo^pOzq�O���P�>5Z����]}�o��H=���Xb�-�ρW���˪�ZyY�:{����]�\B���� �n\|�&��a�YQ�+ �QAq�WfF�q��鵶4	�GD�4�)kiiv�b �37���A9�o/�0��=��>�Y�8�
\�׷�ɗ�a�x�M�]�0c"X���]��!б ���0`�'n*,�M���{�����<b�<���޵Wk�8�:�ۿ�{qկXY�"+bv��^汆���bG�Du��@0��>��!�c�f�����\+��*T�t@�>�2��0�n�j1s�DO�3�HU�w�G$Ġ_����	��}.r;��c$&�{��A+����Rϴ��nJGX��a����g|�ڈ�ԑ��c/����J��x�=�������7\f�<�5��:�|�	{ꩧ\%r��A����Z�G� cGŝ"�3��7Hj1�� )mf!]@����T�o������Zo\"9p�&��3��v���z$U��c�-����y`,QV�#f}ú�Z��u��Z��+�Q�ǒ��K��d�vDn�b�Շ��"����)��]���C�4��U�""8ҐV
�J�՜�'�z������|����Ȗ����D���N��8�rr2uq0/0LF�����!�8,�H�Qd��l�O�fg��v}7�0�;.�)�m[�t]#�!�eA\�tp���Ex�E=f�X?�Y��&)�LQb�3%�#)�������f�R��DDA��e+OJS�ܸgqʁ�4F~%E�|� C	�4����yy�Ĕ判�����]��\ �h��r�h���1��
I ��H�.���'��<g�R���ŕ��/�s��H?�� 'J]�]��|�-�$}}��N��Az�(�c�/h}$��׾�pN��(��P�l"� ��O��Y� 2a���z]���G�ȒWV��A�ΉB�t��o�|��v�M7�yH�l�?������������������ɟ����_��������?���&0ʎ��A|�0A���K�m��@�ĒX$&�!Q�4t6��A���#�K��j4�����	jLl�65�dg�����|[�5�����v��I;|����9z�>e��q�>k����G�ڑ�g���s���8j�_9 ���8�oO��������Gl����������2����H>w洋���l�T$1;��K�����+��ן�ի������;q�=v�֮]��������Α�X�~���ء�倈�5�g��e> s'��"H��	Ӫw�L=%`JI����>WE00���.��X�;2}�_q�߶��������ԧlㆍ�L��w���[XN������Q��Ν/��H�x��:���P�P 8�@g��/����a���o�gڙwBz����,b�c�34|_U�P,�p�_j#��{P�ʱ��^^Z�z` B'�4�p/����D�Ƕ�y.������ ���2����99�߷� p�ÂS$o�*DR��g��0u�?@�����ւh�d�0���D�t�w�8 I������o1\��B�-�H�� ^
 �ӕX���>ho~�]�?{�s����^z�N��0����a.�ds�%�Xrf�{L����EL��x��eiOp���w��]�|�
��ciw���(��ǐ�(��w9�P��:�Ƈ�a0��´9�rT�8G��dX}{��r��ն	\Z����;z��?Wc'���������Sv���?��@��1;|�8z\@|�^9t�?a�N��cg�
h��R��;����*���������s�W\/q�y�����&l�K{����G����+��-7]+�̴:}{R��*�b4Q���H��ыsr$�@���rb�x�N5p+" 8�U.�Ad4���� ���P�3I�#'��X�\\g�}�K_�-ۘb�@"G����з�ہ�|��ͷ����1u/����c48L��!Ӏ��p�$�o1b+�G�)�R��X�L��=sJ}^)��\ý���Ce�}8�D�ñ��w��Cc� �x���%n7�"�����鲫�������/p�e�}"��o�'�NT=��=�ܳ�>辣/?p�p�lP�� ������{�2�mT@��#���r
+\<���=	@������ECy�a$ ":Pއf++�1��M�<�a换�$��4��{=���^y�cF�Q������w�w��"���<#|ȷ�c�W�SG^�^�m�f������؅�xޡ"DѵƛR��\`:H4�� ���u���9�݊�s����\�J����>.R��H��!�^tZ����"N0���rW[A�J+\��
�����U�[��ݳ+�X�z��%K�\e��,���2J�-���X~�l��,[ey��W��r��V[^eye��@�ɲ����s�蝱pd$4
� ������pf=�C1�,�EoOE�/"<@�)D�+���-ӨL��'��_P����O�W���aӅ^( ��I�6T�~��2��k�q����ii�����L�!Fd��F^���	�#0H���rB����V:z����|���H��ի��G\��7G�v�J0����� T�6�NF��lj�*"�t2�3, iQ�XՔ"7H&�nU�"��u�����習x�4����Ģ=��i�1r.����c�z��Vqeo�����~�7�wr����K������z�[��v�w�-;n��۷���,�E�96>�:ol��*օ�'E�V��$7/�u⥥l��9���я�M� ������=�)�uI�"=#V3b�R$���0��f}N(�°:�ں��~�=ﱻ�[�������/�w�ڳ�;&��9Ǜ6_�K�Y��\W��*�ӣԙ�ce�
�-��@؅�c�3�/��@��:� ��mB�~_Ƨ?�)6��m����,)���JYJv���W�31�`��JJ,O�U6g���8k���^E%�_X����s��\#=3���Δ[v�@Z6;7X�a�Hཤ�҆��O��w��uUh� ������Cj���jK�,��ő�s�qG�}���֯[���j��sv�b��L�	����
y����؉�e���"�QBF���{59)MD�9;���"�5g "L\F�A�{KK�z�C�ޟ~���b�)����Z]�ܹ��<��O�b� g尵��|�+C\�V�p87����W/�5k��*]W����˗���*�~�
�e��V��+s7ʨ��Xn�R|��JqTcV���E��a�5z,��i��C�*C5���<�gՋɭ�������<ͧNx���.�	�gz�1@b��͛7���!�e�:�Ū�"�B݆�}��F]� 6o��: Pp\w�u~���Pe��� Gk@��>b�4 ~�Ƈ��y���F��qF����JǞ!I .�Pc��-:V>� .�PC0;�A2����6�w��<�䓾)쿚���p�c���~�D���� gP�e�
.� �,�H[�;%?�r����|��,�8q��#0�l)$6: T���"п���<�9����zb�u��[:��́tZ��aw�%����5M6:+�%-˗g�.��2G%�q���q��I���!`�D6��Q��3�����ظ��	����G�=�$�<*"`��3G�h�r�+�( 鑣g��^tB�p�
5�7_�@�h�2��ۯr e
Ͼ}���Q�����''g���I�[��b�ߎ>�i@�G��B~���5�D��*��)�"�{|�)�"!�p�H�8��*dD0@��IK�8��k��@G��=��c�z����~�8�<�^;s���/��'�\.��6��a�^�Uyܬ���6m\o�6��+7�q�m߶I\�����s�]��v��5Wo��U���ԁe1@�$�ݡ<�5kVز�*�b�*۰~�]u�_G_]�����
�ɠok�X�ll s�M��t���u*�A��f�ިm\FG��е��f,Р�Z9���a�|�Pkj�I���}pH!���d�7T4�f5+�X1�u�V���n�:q�+|�-�C��|��#t�p� ,�e N��( �iUb����3�2j) 	����"��J',��g�"w�@J�F�z�[�b���6ߝ;wڣ�>&ɭŁ��@BC_�y�fV� J8`6;AzB�#\ ����-�T8�8rRZ�},�ӆ۩S��'~�'�r�bׯ�.m�<Ĝj0�z#�/|��5�L�I<�J�^.)좴��O�3X��7�����mbFbuJ��S��*Kg	Sl.��i���eG��c�$:e� �C?.P��L2��e��a��'�����@Y�ĕQ�$�`�%�����{@�U9�D�%����w��Kő�Y�8ر�Щ�gD�jܷ��r�'Y��d5���$
��E��?8��q�~�"q%%�608d'O��h<ať�DVS)�
#95�fE4)��Z|�	�ۯ�N`W�g�,�\"�o�s�p���WYs�G�8�15�M"� 4u�M����� ��9a˿;�]`U  ݧF~ħ�p���y�y�,*�ձ$�X_
�n5�Qc�	F��R0�e��x�BG�w˔'�gMM��W٭��n�N`�сa�8��˪�	�q��U۷�W��I�6����%KpXd7�x��c���J�V��֪���8x���d�|�0��FO�Ξ9�)'��fIϿ��s������������]��ٳ�����wz��w΂gd�I�t�t�̫��uW���D�ܫ��ڮ��%|��,f���� �����FG�`��Z�R#@|^���iYH:�T-����&?ȏ�R�]�],)��oR�T9-��r�1K��8�߾��o�) ���)l��^�i��t��ܔ��/�.�s�a8spU��/Œ� Y6��~�1� G�kg�.�Pq��s}���-�����E�y��K�����p��:�իW9W�Ĺ��$}\,i�L�_9����~;t��&fYq�f��$�3L%��5bߴC"^~N�D�|+U��� 3U��4h�̸D���qK0��vZIS$L:L�ѣ7>ǔ�;9��H������� �r��{��]�l����%Ev��@@Z[^D��iiI��A={��g45�	�T�F������q���D�Ќ5
t�Z.��H�)�N˰��K��	<s򋬠�\bV��8�|qE�Ѱ�mii�w<-mv��1{I�d�}D�Ξ��ee�0�>r�>���y�u������%`.��{w�O<��Nؽo|��C��מ}�)kint��Ν�ۮ�w���s��Z�ٳvZ=����}���C���QX/v����_s�U"�*�Ymee��@�vFU���.;}�Y��-�*�Ԉ8�d�n��:��VT+.*�IhWg�5�:�y�ab�A~'��𬯭s#�@���|ȶm��:u64�%v����.�'NP�$������B��-O"peP
��](�x�l�Wغ��l�8�u뮰%�q�p�H0p}X$t��w��l�u����������}9��\W��J�L�g��u�N2�U�3K��-Ϋz��g�董?�88g�P0�����G��x�=�G�G�w���[4�R� ��(�"������t�:{fp���H��� �?�@�@$�� Q������is �����mvX��,��^Ƨ1L���`�%�ZYn��\Rn�W���ն��Җ	���1�g�\3-O=�28�qG���h�|3�6l�*�f^'s��
�����le���
Z�Z���n?��S�}=o��&UH�*��Ν�ѻ��r���T ���!�ɗS�9�q����aMM-v��Ab]�M
�S���R��-���)Q|\��T�u�Yg��ut�)Nٮ^�Y�5�t؉3�l�t��X�8��e+�����ڶ�W	�3D�f�<��w\:8&E��eڑ��=��z�o�[v�j������\b*��^���聙#ȕ�����f�:�3���{�5�@"� �Ԑ�؄��|���lGx��qo����t8�3�u��p��:OX"8��e 8Q8�$��u�ã��C��`MWg��w�}���������}jΒ%K�Y�	�pg4&�9މ�s��-j߾}�`�Ӓ�(6�fh��p�˗/s���� � �J�)���	h���2%TLM��U�QI0$P����>��/�]��״��$Ѯ������)��d@X5���x=WS��N ��ԑ���Yu��755yYqe���F��Ĝmt��Q�@��zf@�:NT`#q�Z�-z�m �QSc��b.!��P�W�H�`����&�i�%��2%dvfҦ%jg$L��ťv���v��5�|�IN��d|�7�"�%W`��<Eɜ�L)7���͸���rD!E��&ԝ�� H�:G*�J�s:�����/�GU�Raa����V��#����Ev��kh�s�VR^ik�m�ə�V����)o�C��܎���0j꭫g�z�G��W=� A@86mv���ں��hZ����S`8#�ePD�(�E�'<Wk�O��s��ly���ű�:�r�1��Ѓ����R�)V����[n�믻^ �jǎ�~Id�6��(nc�UK�K*���k��ڮc��[܍���}˕[��zW#�!��o�������o��7I�,���)6,k�	�ƃ;F[\Y!1r����p,�[��s�`��0���dr�o��ڗ��e���<���b�O�s� ����kw�u���\�Q����XA���
� "�^�
T"G����P�G�q� �4\���u�(�V)�`72�D8�e�
�q�G,{�"R�9H�6�Lu�rr";,��?�@����F�gg���	��E�}��a[�nq���'����:�p�9H�;e3I�$8���g7��F���E��F�}0�y�
˗˟�|��,G�pE���>�~b�,>��	�
��b@�9ЯE+�H1`ys�h9���w��;����q���N�b��*���d�"q�k�Uڕ��ZuQ�Mu[k�Ik�?gý6>�o���T���>M�%z��l>��*�g�
�7^�s�/A�s�X%.�@:* E��6dƨ^ŭ	Hw���LX��iA���ı����/�+"��{�H�[63	��O���B��'�5uv��I;#n���צM�^b��'.nd|چƧ�wp�ݧ-�F���PS�ع'��F�Y�����XR�L\�2כB��Q&9?��3V�^bg#\��dD)�t��m�R���z�H��E��T_��J�����գ�+ۗU-^"�f��]�^��[�c=��D]��J�K]�UXX��������.��9��V>	��-
w�h�b��=��@������*�Q3hA8tz���EV�h)[�@1S`���჈��>/���$pgz=���r� v3p��),3��ϧ�2b��6ɗ��#.D|F�Y���x�?Ɍ8<�8V>lޱv�Z[&Z���� �lN9�d	(�ޠ����,v��iGp�^1�hSo�����Nv{���D�}�u��B=QV@f��k��k.4G'��+��.p���*-LbY-�A�P�W����΃�w��%mtD����{9:]�\v Uy@K�׭_ﳋ�̫��oV�و^��rB�}�
!�]�SlU�"۸j���u����4�Z�̸��f�hn~A�z�|��ϲL�����<�ʞU�r�(;9ǠODi(�eBs��l��^ ڗ*�Bx���Ў�}�����&r���?���F�텝/�#8��L�$��?Ww�u�]���fum��8�{P ���N4�Ƨ�6�+I@g�ل�z�4))Mib-5ǭ0�/KĞ������I��
�1�htN�~��n�
�d�K�yP���ƻ}�75-�N�<o�^�c�Y��p��Νs�#�Li�NRCsK�8��w�J�Щk��xO:�����*��q<���lvڮ]{]���9���ټ�����^V,�?l����}�ŝ��;�%���Q�����uYL�@��t��E�I)o�&���ږ-[-Q��@̳�>�p�s���Eғh�BX���%"9`G��+Ζ���������f�:c�ӋN�<�m���(�j�a�2Y�	/{ ��(���-޳i
�B��t뭷8X.�}~�S���\��N�%k���S��|w}�	]-��j ����6%�/���� ���3�ޥH��� ��9�銃({�4%/'�W7�H)8p ��ihNP�颴EG�0�I���߯=��}��-5���+J��d��U�H����`�gO�f����K���@Ǵ(�Q%	��i����.����k�X��;�Ɩ�v6��H���F�T^�mug�`O�}�_��6�_��oK41���/<j����n��zp�^+)ʳ������8g��͇�muj�Y���;t�� j�ŕ�֙c�gf,Cet����N�ix�Z�����q�x�S���'��g��1�7`ij8��Ɋ0��?#�ɧ�F��9����(�:C��)v��p�b�y��}�{m�M^E�w�f����9&6rF/G�bfBnN��`�&��,+J$�{#�`�$�g��A�pW�s��9W�Jj�	����5����?�t�
X�|�~����������&u��"�YaBG�,X]^#�U��N��d�z����~۽{����|̮��:K����������m�r��0�IR~p}S��b��BFO���s7��|
�f@n�{W���3@�'���z��}�[�j��s�s�p�d����p��t841/'ϲ�.�Cn�&��������P�w�ޮ�j�}�������D?��x~V	���+B� �����t!��.���Q�nv*c#c��C�}��33d�9,_����� ���c�=f_��},�K_��:}6Z_��0�y �^0��_������c�g@��q U�0�wÍ7�I%O��<;6�q%��^��_L���S�������]��8���4���J+m�}��z�u��I(���/� !@(IH�j�{��������5E3�F��yޫY�lH²�}�:�W3s�ν�{�s��=oI����P]Y���L����h�l�"�8/'��*�/&��Rx��=���d(��V�e~�70Jf���n*A̕��¯MG�NQ���@V�m��u���b�^R�:��"��|�;��S��+v�{)��'C��+_�<6m\h�`�N��yGl
6P;�lWeh���iu�]&����~�����G_Dg�x����S�K� T�1�	n�{5ӆCH"�5�bt�[6�!���N⑮c�%;�؇��g�cl=���t=����g�́��9�HM�rTd�
��eG�Q�������9�leӧ>��Q��I�c�7tK�& 3S�&��R}�&2��@RQ;�Q\HX�^/7;M5p����oc��ط{���u`;+���*r���aݚ�u�
T,�������ٳ���}����~����6�����g[�Y��LO�M�OlU�N������5-Z����~UR�ذ�U��l�7*���.�lٌ���L�n���أ���g�2p�B����IF��*�=/���r㦍x�;�i�/\��~�3�ڽ��5�V��O�i8���bں?�Lk�Ϋ�{�{'.j�̮��J��K�U����_��cl�e����s���^9t�H�ŷ]�v�G�7�h1dUr�s6�W��UE��"��ƈ��Ƃ�E�L�K�s���8�x�bQ�_]w�w�F�!��6t���ŀp^IJ�30EQ���I��������{]FU!�	�)ure��E�����8�УM�Aќ]��-ŵ����ѡ��}x聻�,6��J�>t�,v�9��R��-ݫB�Ż��)��|��8�]�H���$�md���OnnǸϣHPI��󢶩�Xr�#��(Ց��޳iٙݬ�l�R�{�w��A�[�����m(+�CaQ@�����8���m��z�����䳛 7@ȿ��(C
=��#��na���d�!+�u�٧fd�~O�B��RfOni�H�-�ﳐ�!��L�N���dMe�$�\�P���=�����D�#���T��<>�efv�t���w��J�N$6��BNvjj.k֠��Խ\�r�k��K
��X*���KLkm�0��\�"y��A[MN� f�IN,Eb��P��F&⫋>G�i`JWj'PMJI���A
x�P%�nf��vVp�K�v$���:@+�ÜLeЮE�u���}�~�a�Ks^|qv���u�BIq����h#Aޏ�;�(F���A�u����������j�I��kr�4$!k��I&�+�����I������8�~w�S�D~��7=5=g[�f��y�¶y�*��E��߫AT�
u�t��Tl-#-�|�>>��߇���Q�v؟B�i���Z��;�����prccFۢ��eKP\R�ܼv�4[!�i'��yf;����"�$���e|��/;ɚ�zv�.��u����N�(��Tn{A��<�f���
�d$d�d]`fB�]��e�r�!�H?:il81�py��Ȥu�$�n|�P����٧r�g焽���<I�����،�����foŀ'�}Hg9Ȏ(���������~!v��<� *�����Z�7�\�j��'��]�:MI�}ھ���0���!�4��������(�/F|ܧ�P|N�|�w�9���c8���q��9-�6>�S�"�����ױ@Ԫ����U�FA�������f�/�y�i�) �҂��G"�����X
�l8E�>�ҡs㠋+�@F�d�V��_�V�5V<�o�ۦz���&����@����w��ݖ'K�t��}��Ac��n�ͷp�&r�8�G�ϡWA�6�1��&��5�e�(�	-J9v��9�إ��7vTI�bi���R��F�T�8���,I�e����;`D�\6!E�G�ME��a�׹�9rS=����KQ��'�6M|�����r���t��u�d��d�XT]���l�v�`f܏�*ĳ�464q��ɚҬ�����l y���TtN)���+l��$�9`�z���'9���Z8�H��}O��w�2R=��#��;��9�+��}}]h�WB��8i^Agm;��4�s�.XP�V��h�|����&555�~���38p�<��'���K��&�Qj�C������T�V�'M(�h�>��C�i���UI��9��f���c���^v�Z�QJh�sljnŷ��ctt!���,d�/�"M6�1%f��Sa��u�Iv^nZ@P;*��mS9�������L�l��I<�2����98�,����Plu 5�hHP�
��k��͠����=:t}U�A��W�/�w��j`K7\T\����X�v�YWhe[��T�X8}�'$h��tjI":�^�:5��^�)�\�S�P�"zS-HIW�WlP��eQ��o�kAR�N��"���KK�l�rK-���[�Q��@�Y�s:q"��?����`ǎ�(͌����+]�R�8+�
{� ��z��\y���r9�ҽ�0���|�s;1%��c�)�U*���>Ug�K6���A�tf��5�����q�@�jk��,��u�%��^Ϙ�W�eD�Vu�s��{��q��	421��\��.
��h���x~���U���6aqU!��o_6�ZOz5�Kd���LQ-�Т���Y��YO��Ըt������<���.�t�6ӏ��R�x��O�!+=~VGڃ���?`٢*ި�#%	���{��?}+W�5�=5Ń��z�f�� Gx��QvTͤ� ����s��(N4('����EL=d�Z��+o%�rc��+�5ʨ-R�s��5,ZK�(>fI�d����-5�QQ���x�G��,�8����CB3�D;E_�$b���n�,FrJ�+��{`Y'SV${�1�$P�OUϢ��ΡM_�{37#��ë�^O��Ǽ,��M��Ų]'Ӕ���/�$%E$ٙihm�GC�E|�ÿ�m7mAkK�� [6���y�
��'�{��nq����[��-������m������/:ZT�~T�b[�<�-�����>�o�/�^t��W�=�@E��>s��%��r��5븪�*�X�ʞ��K8�Ů�gԷ���F�9|ǎ�$�;�`"��K�� X�~��Uw�_�i�Ķ� ֏f7}�Ģ\Tr�{޹c����V�'tb��f���6$�F��}��I��*�������n&g
p~��S]��\ԎN[:E_���f�omv��E�N�W�u�Y&p,:}� ��,5��WU��W0R���2Ҍ�,,ZP΁����v�y������%~s��Fq�0�"Aku ��8�Β��k"��0(���KQ��ٍ�7���	�G�05�0Rǳ�aj�������eQ��z��٣�p�>�����6
���L�2��D<V����A��j����d�V���"hu`�
r�	�I(<��E�'�#��io���W�u_�d(�= �#*r��\ʔ)�Dd]�N�@aQ�]OI�Ўx�<p�c����/���d�n�9�G��z�M��;>��"��)^'�g��S�U��e��I@a�t�6����Y�c��=q�7��,\a:�l�ׯBq^�#�M@��~��E�2��:G�n-��eQ�HlP ��Kr��兀M:l�����t�׫���v��gE���Tmyv��|V�Fbwb�Z���pee��G�_ʻHv����z?vgΞ���N�6]��>G)���U�Vc���F\d+��5-�K�@�`�b�ؔ�NJ4'[b��&9����὇-����n6�Hy7)��/�,�Sґ�WMR���y������dff�g�H��w��U�Pb�j��.��u�%��oR�i�ppF�8'K�b%KǬ�fq���F��?6�ǟ>�g_|	��W㾻nDey6.�>����(�.@�;�|�]ll-�N��͓�J�3�$��b��mƔ�X�t%����������	[�q�'s��S,�!=5Yi�ho$#����d���I��H�a���G���	<�f�|n:����G�����@͊��=���� <��$��W<���W��O���3-��|<0�Nb�Y�Ɉ��2�Vh0E��x1=�'{��3'�fe���mHt;���lQ�P�5(hZ�sLIFP���(�7������oY����d�Ć�B���)W���>g�ξ�K������:�3�u�B�9fSbW
�b��D,56�lԎ�U��y�~�@.))���G�"���}�o�|�Bػ��g����\`�k]�����C��Tʏ�?����ޚ�G�>,\�����mj=��Q�I�\���`D�bnj� k��?Hu�}6��8�^��eI�f&mt&0�AD X��cbq2���ICB�tHa�C&B;n�3f,p˾��W�]y�	�!@ݣ2)�;Jj(����꠺:V�|����ʦ�ӱP����Mb��w�ۀ�G?����
��:u�*ǽ��ة�K��SX���$��dYݟ�9���X�~������9�:��+���Jї�����jL�V�W�VW�3�5���X��E�8�� 6��_�#�h���+8r+��H++K�p��vw�qF!;#�I�X� b$��ú�O�dzN�LcL|�X�����N�6���N��O�D�ZLIH����-!#�=�1���{Ɇ�y#e���q�r��75��!�����ؾ}+22��eޓ�č�����{��' -�C��--��d����������E[�b����l�?J��A*1NE���Ì�!�c��ό�0��`o'������� YA5� �Ջ�tiH,�o����ee%悹t�b�]+��5 z�[��[��������)�$y$A��a���݊��YT���TG�=�)���Yb�V��.e�B�<-�@R�슊/���-�)O�X2Py�)^��'_��l� �(M�"��-o~���̡��]�T%��[4�h�8RQ��A ����8*��e���t�N�����{7�_g�����d�\��S��$��:�&C��/6�qg:�����c��N�_ *�W����&�)�SPf��I)H��$�@V^U�E�H� *=�&�	@���P�^�c�0v���}^������)����8���>��&����A^Z���
Du�Z� �Hm��c_�&T�E	ٟJ�����a>�Oa,��<����E_�������;��	IG�^�7dr�M����_�*� R�X.^nBKG.�)�R9����f�$i)�آ����eCi6W�$�k�S�	��IG)cW��{ !)g�� 1� ��U��J�.��-���[�� 2��p݌�aמcdɲ���j(�{�����4��c<Jnz���4����dP-f�d'�pV�epl���v�a�Q����1���� �g���s��"p�>�3'pO	<G�@��(�f�AlZ�
�W-��(�N&f�
�X�qY�D6�	��X||��tk�h�$����G�v�ߋ��)Q���u��
T���-��ԝSdS�5�l�n��@1:��#�(A��o5��wnwE,%��~�)�IB�g'9���;�07���n';��{��3JFGk3��dݴ�p��=�C��-J<�DV,r߾}\ZU�P���(,���dCfx�J�Y���mC�kk���mQ��<^a��f�I�����4%�����M␝�t�WoR�tw)�G���614�������:�ִ����bK!�c�`o#���F�Ոu��2������ '� �Z�~�������A�Q� t@�@��c<�����W>���/@���E���I<�8��* ���K҄!ӭ���=���C���$S=�^�� ��~9��vy���Yi�W����+�1�Y�������D{	��:��h<��a����2�b�|�\9�h�?�ݍm�WP��|�5�t��&*^���0!d�)������b=;�H 'N_�'5����yB�xZ�������1��?���c~y	����������]<��C8v� E�D|�+_���b����f�ڵ�/�8"�"1b�K��!�H7��� }d��=�ٷ7߲]�]x�٧9t#�3�l+e��hQS|�X#�h�r�AKc�V���q�z��ky��R\��5x�Fމ�����Ǜ��@o�;����৏����`�|�Uo�>Ĳc&P�'�D<[y'ԉ(Y�F�:�:�c���	 Ċ�i,f)?K��W|Y4�%u�ȠPҦ��$�~���{���X����ob��58}��	�y	�U��W4q����vbQ
��Kk�y��o����3�$�l7�]�{��C�����cu.��RfO�>��6Y^�בI��o-fi>Q���\B=w+�-����k�%�>]�E�C畮�Y0�![�5��9���N&/&-�h�]%
i�e�u��svn���y;�8�U�u��s����N���|'�ط��Q
6����șx�������l�|N�
���U@z��aK﬌O>�ْʇ��faQEf+cE_���fQ�^�����WWt��1f�P]]E)Zj���_��r�Fc������GMFZQU��+*Q�����:4�����T��CE|
5��
���b2���I
l�/��mx���^2���^Էt�o�bR;%d�;�c>ē5�g%��<�m@�-Hy=$N|������?q�=�����PJ��~�s����t��o��ǟ01G��p�"�&����
� �;5_OO��/��n͊�����(n�~+��8����q��q��I)��Rn������|�ɥ��J���<D��l�2�k)Ґ�VduM[d�haA� ԉ��4����7[�&OR
�������BA����"d�9� Se?UpfR@kMb��YH�j~�3����$�:+��q�:�&�$-*.��,k��Hu����6����Ly�g�,�p�"��M�h �R<K14^9h\�b��FⰞ��4�/]�W��Uk�
�|��!S���T2������D/}���;�K�+�1�������s qKOϴ6��W��������;�P>W�&=�H��3�9���ؓ�*�*� P~�����&��RU�=:�@� *
�h���r�d.39ſЫ��&�H]�F�P��b����{����+���Q��r���/� K�A0�W�K�U��J���?F�~��aՕ��i�}������}=)��h���⣜!���1N�~�:\Yl"�E��{� �?�(O2��QR���EHO�FoC��)�F�����OJ��ꎋ��Z�pl �����Qp�DKG/[;0�M6j�Ed�	�(:�g��?��YF:��c|��_�w��c�z�m8{�8�.��/|�(/����S|����R>�X������-�:���+����Tz� �M��O��ѓ)J������N�:���N������V�r����%f&�E�n�hCEB}��Mo�g�]�5��)V�]Q���$]�>�A|��干9��_��ߡ�lI[cS�46lX�M�
�m�&&�mE�ҧ(��L�İ��_\,K�L��d��Z������|��e6z�>��fw��lU���Ɖ�H1'�f�C����3d��X'镢�1�g1�����Jo����SOYd{9�hb�7�V�eW��Zb�]MTRU(١"��k���&��'�R���
����
J�A4r��*��u�������l�b�bNқV̫�q'���?u���	����� ]��O��$.*;ꃇY�%��lQ6�f���b>?�`7��Q�U�/���5F�ҝ�:F�����Q�:� ����I8RI��@�v�:�����k)��+����|�v�����%@j���)�	Tʊ+HDY~����U�h4�����ĥFĦd8�g
�r�����^�ϝ|3�9y�Mס���4�
���œ���Sd���n���a���(cwٞ⇺��~�!ҚsG~!���~������ƛp��	lܸ
������0_�ۿEsc#~�����%�+NdY�L�ג~J����/_`�O)��E���6�{��K�s�� i��F��9����إy����_���� ��cFb�#�<b����5�Lv¦�&|�����O?mf8
�q��������N��羈�<�(�1�����i�Sw�y-�2 ����d�8;y�1�_���?���kU��<���b�����n�)�����w�>�6`� 	��I�/��鱣G�H�M�T4 �U��+�6��Q;�	���t�
�{�
`"�5�d�6�&Z�p-	����5s7�W_��E[G'��̗p�^�d���P�"�T����+����y�z�Y�PՎ������K�Ϊ�*�<݃�[��䯯�����O@��54����.��p̦��ʙCV��$P���#�HN����&c�{��1���Qw���f�Nܣ~�xH�U\��4�l�|�0��7m�JP�g�O�O�,�ZF���1���߾.��k>'�M�.$��^SgEq��U��
;ґ�j���Gt�eb:v��0���� �Afj:J�
��IV���������fk[;Y��E8�̤�F��Fwߐ��D�r�n��Ģ,�9qrB�:Mv�������,$`�R��=�Q[�H�)�u�Q]U�-��s`$���#(��!x)�O2;�����LPƙӧ�i��:�xm�M���!#%yd�9�Ɉwij	�{���x�a����#X�h!
)w�)�QT�O�������=fu�S ���Z������o�s�v�Kƿ[6o&�L�����+J��ğ5�W���>~��ߓ9v������=��{v���'��9??K��a)H:��'�s�9�"�D"�M%�5 S51t�T%g�s�<�
P|�8A��0��:�߿�k�*��r����^�b'
1&��t��Ճ�7[�[����l`ٷĒJ�8�i��~O`��"HP�zFK�e��G&�W�\�@+P���b���.��Q6A6^��D�o���t���n�����f�5��!��>��d�t\;5�%=�dO�4 �$�Ȧ�:�|��M���'�_ZZ��&W�,�1�Wmf�?k+,?s�������8�	Ikz�M���!RG��*K��Jv��%a۶m6.dSj��%��nS��_�V�[~����Y^pS�lIgJ���L�*���ZR5��OƠ���=��! D�9#���@BeSQ�T�+h�fO�k"�')9��؃o ��mhi�̡�*�S=bŁ����փvqK�8@�U�7�
H'H�v�9��5Ypc��*���Mk�艷����,���4zp���]IǺ�;)֥�7�f"T_W�N��2���r�k�>!��b��;�1��|�����w�f_�D�j�e[4��ut� �����j���?��uZu�#dl�?�����λLu��N;w�d�$��h�M7#?'gO��޽{��)��[�l�ߺ��(�L��C��>h"���47����O���=�K;w����s�>��	~?���q���A,F��l��Պ���:�ٕ�j��]鉗/[f�
�M�eJ�뮻��,���EU�,Eُ��׫X�'�8li��x���ا�D�F���n��D�D�F�=�X0�M�V����e���*�2�J�1}!�k�Ɠ��k�M������)�4�c������d 5�D{���إIAj�趶����IOF�
�W/���G��ڌ��\�p�/�'�l�8�~�g�.JF���q�2/$m�.���#<�Dh�@'�m���L�$�;�؁.JZ���n��j�i"֦�~�&�$&}�$�)�Ì& �pD�ޯQ�i:o�G��^����"\��D����~�:P�דuD��`�sH�/Ab6�h���cH M.LIC	;PA#'K�=���Fc���k�����o!����y|�Uر���Jp�Rlsꃇ�������Gy-/~JѾ���U$��w�C��>�e<�܋����������ȇ��g���X�x!��[@PG����{l�`Z�x�e��8q����+�˭Ì��5��́�z/J`���",�=ihj�A��8n��A�t��{���8K6��K�y����c횵�W��>2O�W�O}�uX�A����5�����V���(*��?��?��������?�{x�!�w%t}��E��҅��T!�$~K� ��v�:���1��,hI�&=�@@���� �ߧ��@\F�r��ѵ��Y\�I* ��m���I�m)�Ů�(��S�g�O\��ʲ?��l K���Cz>}%?o�3v���Ģ��5�O,5�CB�>�,-'0��O������JN�@n~
K�LW�(ZG�_8�x}1 ;��E�g4!	�496SB�j��P$��/��e�$� �u�y�u�h���{/�˳~ �"}��o�b��ħE&'��TW��&�i���:ΐ`D[�M���Yז"1X�c��i ������(��I� ����J}J�#�2gҽ�����/��.��S���Hr��XԊ�+m.�F�'2�B�W)�@��#�c�������C�41��ʙ0�8C�H�'�p5S����1�ef��N�N�W��F����S�c"�<�X��{�&�����������H���3G���o���0��Dw��a� ��/�-�z��߰���[�����.���W�j���o��陬���A�'1L��|��R���RCm-�� �+�U�A{�L��A��0�f�$w�����3�^xR�p�}����©35��o� ��l�[������z�����Ϣ�=r����ZҾ���/\��>
���ގ-7܈?��?#���}�o�o���+��n�q�ٍ64��⹋(-*�⅋8�:���!�&�$�EǾ��ا�]Z�U�ܕ�L�B"FZhB�32��O�"�G�
H�2s)��+�����Q����f�.��,^Y��Q�K_�������~�֞�l��βN��[\m��J���4�.Z�7��
,��'�&����0��v5	�?�u1S���D�g#+����gglNϞ��>�{�~�G}W{4������̺M�2U�~�_�~�^g���gk5�rΩ��O�O\f��\�����5��z�/���u�]`zu��\�����'E���g�g"��{M �04�(݋bh�-�Z^�3�}��	љ��dc�s���:i�'8���F�'��~���ű�m�I���2˱�R���h�X�4#�����R����4��'ƣ��a�[��?� ���H�w�t�N��������H���/��U���#����������J�����做FE��+io���z�/�53�Ρ,S�q�OGK'�icݜb�;@Rzn��^�K"��E��O�{����7�����n���� �Jӑ���=~��G-��ȨO?��E�9��oߎ����QZ������w_�됀��������8w��;O\

ɂƃ�F�sP� �Q�����Α����ԑ"z:=j��D^�x���fUXPhVj��.�a��$$i���PcW��	�����w�X�f%��3�S�U���g�F-���gܿ�^�Vj/��d���6�CĺԦ�J�#}�k��Qd��)������*�j�K^���)3�B��Jr����� ����~�b�;��sj����}Dw�ZE�7�E�P(MB��t.�3��lO�2ﺖE� s7�i��G�y��P�v��$�*�5����H��� �܄��L��H��Vn9H��M�FQ�51�"�:��y�G��e
�7:���Y���M��+`���J@*��tO��/�@e�����
H?��_Ó�<�u�Cd�o����/�_�җ����o�N�7�ߎ�gH5�H��KL�x6��m@χ:N��AB��@*�v�X=GϦ�q�\	� #s�a�ֻ���CG��ŗ��]�\f��?�i�z�<W�a���VW�h�;j��}H��t���V�?��O����7����w4��y%X�N����Pw��"jJ:�X�Z7�Q�MQ����Qtߕ묞:`�}�"��`����l��0!�Qi��'r�cC� ݱ��O_.���Gq��w�g��i�["uD|}��H��]���t�~��j�r Dm���6�>G=�s�M#�T����y�iw8����p�9���e��-B�k
�m�ɾ���V�����.y�+߿VyU���O�f�������0�Z��1�ͷN�%��n�Ŝ�֬]Gv����^l
�5l�E�l�B7͊��(����%�)ʤ��e�� 53)�H��� �w�݀f$=t�|��3�])z|ε��}Eg�G�,���E�4�K��J�	8f�:5)�.�<�d������KS �յ�Çl�=��t�:���ٓ�\�y29Q���ʦDiw|,2�S�t�����>�~��غ�fs����m�����<��[l����֠HJL"��j����5Vo"P�aϾc��o�Ͼ�]�^��08:��d,fb�)vj<&��8|vN)���	ʅ�<$�� !Q�S�=�����K�3
PX<E��$)�	'�INf���$��]���B������y�VZV�%KVP���2�)���jX j=�]���n&�ڦ�|��T"�@����u�R��"E,�LKO�n:Dgs�"�#��Ч�m՝`i�,� ^D�$)� �g��{'0�>�j����_Vt�k݋t�&�h�m�j�kn��_g3��+��&e�L�!;Ts��]����C��ϳ�6�>҉Yj��my�颢�*��37	؝��@���E��I� ��1���
"��d�bqQ.>��6EwN���η��s�H'Ѝs��s
�+o��^G\=�q�C:;gr��tt:@3�h��n��\�R�em���"���ELK���O]|U�[nQqW�s̘���/wJ��Ɣ�y�B������\�Sy�ԞJ�v3����%%���h�%O�O��KJ�F٬i2����+��]���|�/��E�PZ�Զ��P^��U��/GfN1'�|$��x&&g#� �!�&x2��}h�LG}a�����{��o`��^�8��!�(�}^���a47wR|٦����DN-n)z�D`�y���� E6vB=���k\gAU����3� ��X������E��A��m�P��+��9lR��X�d�!F�sɅU:J�+x2�(;���@���?v��*W����H���-ھ��x���f�U��k��?�.Ц�ԍ^�ⴤsm���:*.��"�4~�pz�lqW���'˝|Q��a�2�K�r��ư1�({P�`p��X�� ���h�iH���,v=^Cî��v]禍�^U�Ll���IX��Qf�g��)f�kni5�0�;!���#s�iX��,�ƹ	d.��g}�˛��X��rw��$�(�啖�D^Yr-��)�y=-:��V���cf��� %9�H��6��vT�v�j��i�|��)�<i�58 h�1�Ĕlc��1��?��$��3��(�mjD��_4
J%�}�
��.�t%��cF	���cb���4�$k�������x��}J����j�Z��/=���kE��^ԗ�dV7%u��^�@��O�ٱ!q����6~�p��#!]af���ΜM��x�	T�{���n7Ɛy�ƞl.%I��}�ө�kg<�*�옿�����EV��9��SK�[������;����G��MR���V�$�P��u���6W�A�U�u�!j&Fs��ة<,��lS�ءf�1y��m�O@�i�}@v�ܮ�j'�Ճ�ݶÊ��.o^�����1�[n�g�C�\�l9�ߏ�A�=wg�y��ӏ��V��w���I��b� ���wr��%qK�CBrR
�������\�C���x�UTc�ud��l��:x���:���?!��Q�K{EKK��x� R/�NR� ����	CfD`������U@&������(!����=Ql]Ab"�N����T��_뷲{�w��*
�t���Q��t.��K���(�J��J���ݓ����S��$Jba���ы�1�
�j۫��n��=,�s�.��R@!�� �c�~i���Lg*��2F���l����&�|o+�|���z�c�y�X�S���~Y�W�gݍ)F66��+���ߩ����m��v��������ݟ3��#Yw�4�P����^��\5��N��}���fk��U#]\�ɍM�tJ�be�k��\s�r�;OM�����~do_~}U�%��h?;���_��G��DK[;�4��?�5u�bM=�x�y|��	������]�p�|N������̅�8ۀS�p�B�]nÅ�.\����^�6������ǣ�������S/������ ^ܱ_����K_�
�?q���������)��N4xe��kaŴj�٪���o^�<T��@��U"����($���+��&%uf�1��ڄm1.K
RE��2�9���(u`�S��~ֳ����NP�f�`�X�Pfo�Ū�E[�WlT�tư����Sy,�oP�0b#o�"��lQ��{n��k=�����u�>��l50�+��M�g��N�M����{����r="�R���T�S׻�k�fu�%�/+�a�W6��g��m:�]7���li�бW�6�_��<7���Qu�?�����=�8]UT_��)1�a����Mh% E�E�5�4�_3X
���Y��^��j@c�ܡ�g�9��l�#�J����	�ht�4�� w�~+�A[����<ݮ�G����pV��
r�~�*�$ɋʏ'�|�W��������G�`aQV�]�Ԍl������c���Z�{{�p��q=q-�=�khCcK'٫�@܆���я�	��/�k���E{gΞ���{�����+,��U�QLq_LT:PE�#Qvϓ'���G��MF���s��3s�`��Ch��"(�Y'T<�� ����b�d0���9�������NDe�!��AW����l�d4q9I<�O����11J=O0�-(��d�u�y��EA���d*�<Dz����M7mFnN&�ۚ9h���z��s��Ry�0b�>�~�_��rUofq��	������o�_g�w��?�����|����Y<�W��P�W^u!g�+���ZۯPt�m<����1ײH=����s�+�_G:�/�7>-��\S�����b1�`ϝ�~xeV�S�y�!��(�(��m��}d����Fv;�U"�s��t�*��Ħ��l{�^�t��DZM�����cv{2ux�γ����/�_��ۨklAN~�s-U�'�.��e+���O�~
��$S2��S���lL�$c|&��|�<9���g���x�B1(,]�kn@VN)���p�5��dl3�(K�MJYq��)�q��)446X<�o~��η����ZdggY ���L�(E�~R�3�Ѭ�Nt�D3�8=�i�٤�����icfQSA��D��HG<6�,�-w]�|��(*�����<J��_����Iܑ�J4�f<�R�ߵR,���&B9����B�h�Q-FG����#&'˃��i��E��+��{��/�+c痝MǼ֦���ڦ�Ƣs�6���]"�nE��^�O� ��Dp$��V����Z�����r�?>MFڌ��a����#uD�Rc���Ћ"8Y%��8���	D�{���{c��ڧcUa2,���G�Ow[�s�q��m�d������q�R-�9�(خ�o�q3I���&�ĉSػo?N�9G�j@}C����� .�Ԓ5v����|��tuuY�'�o��9M�E_ H6:Lvڅ��~tt�"06�s���%X-�����c\�7��ϟ6�d��;v�(?�7��.�����1o�6:VNw�}'

s��Q�OV���ź���Ld��9Fp�A�¹�QFS2����t�LTAH/S�!e�@S�죧��bRiS(h!��T���33E9;�����y�0'�i�}C|�M��Xn0�����O�8f���ʶ�e��qHg[���Gb���j=��_�sϾ�7��ȟ+����VI��SEß VxLbL�Ȱ�j��q���)�$O� ��4�}p�I�@�Ah�(������T9�0�;`�> #��:@�S���VV��ˣDD��iW;���R�qʟ�q���:}El��e��]wnGV���5� �ő��<TVVY6QS(�,hk��)�{S�O:��T�W�RЂL��ZZ쵸T�c��j�Z�ͫ4p�t��}��J� ���
�Rl����_z/�P��O:Fy�ȖP�L�&��|lٲ���Qu40���݉��!��吡���2�W�{1�{�����@�C�a�׋ _��A�a���=٢������+7�����	�3�w�V�K05UA�K>���z����Dw�[5����m[���(//!��*�T�J�3u��:�\�+��"��b�#�J���Aɪ��\����$�f� �%������w������,��?H梕X����	,"�|IRDtXWOp���]#%�H����J��IV�K���M����'��䁝X��_��_����
�j-��]��~�o���������<�*x�W����Q�����Ĥ>��ՐZ��)OT���~<��3ر�%3�X�d��^�|9r�rq���S~�T+N��Qhǋ;��ނ?��s��c[�ޣ���b��@!
ۦ@�2�WD�)���+�IJ@SW ��̗�P��ze�>�d�i�f�t_DvZ�󊐜�
O|��e�"{�̹�
�at]������BdS�4C�e�%�����`���c�2�Ҫ�����"h)�������m���|��m-l'����,D�A̕�r��,Y�R�X�⚢�-Y����S~�@*�>��/itB2|�i7�AMMm��Ra���,UI�Wx������bd|�•V� ����x���wb�B�_eE�<��R��������ō7݌������ן��s�k\dyZ���@�	�'��Q���:7�=�
���	��_�� ��x�;�%D3  ��IDATD�R��:�,���t�+j&������w��C��_�b��Y,|n-�a���W�D'��ب�c��Xw,j�|���}]�~����V��I�җQ��[n؊��"/�Ѐt&��J��A�h��f���?fT-`������"F�BS m@��\���+��v��$�Z���/0��pi������ĺuk9�'��t��y�o������̕�r݋�y��TN����,�ӗ�So�w}��W��)#"ڕ��`��l�T��D�+�6j�^&��?W�ao�$zc��)�GGz��+G�;�'��{� ��ơÇ(
w�wR!( ��
 ��<��#�;��>]�@?:�k36�$0/Fzz,Y�Z[z��23��|Y5Em ��-
)I.,ZP���,݂"0���,b����[@��6Q��&�M䃕��s���������$�#�c���]����ַ�	�<� 6�_M��
f-]��(PJwOz)�w������@o7F)��}ve�AZR"�2��O���'�($�V�V��p�4._8�������8y�ߟE[K+�{��b��3Q����,2�$(OWL�&��ҥ��\��Eb��Ȅ�n��eP���+:R��#�b�(b�"�M()1����H?�)!���l^!|/ݨ�.0u��D݈y� �em�bAM!D�N[l���nE���T(Cl��G-��r1	\Z�<�A�x{z:ͯ����b.��ԣ���"��x)�N@�e������3� Ο=��{��.
�x�[QX��رs�����U��
��h����j�2d��F�M�bמ�X�tY��:NB&e�/C��+�'�e-�;>ՆE֎z�#�q���������哉�qΌ���2V,��#o�����,�h�_��]/���ᣇp��i�>y
'�9��:���h�'��� �DuR5(O���D�ʚ(i���56�s��">�*�0�s�vRE�����(TFخJ6(�ǔD3���\�+׹8ء�
?�
h^XTl��/�e�?�O�E�b�'ԡ�?���|'�\jEB�D�8�$ҋ�LO;��tI�q�'96�Y"�Xb�� i<	4�! U��6��0q�Rbx��A?2�]8��Yl\����#?;S"�A���Ǿ�ǟz�n��t�Z�ӂKp� ̛Q��X�@�|*�t���8�^S�̕�LzQ8�QXﶦf�������|��HLJ���6��׿�Ǟx���Ľ�e�<q��}�1�ş��}�u����اPZE&��c�OA���Ťx�
{�h�O�=��m��䓯 �m��1�@昉��~L�F��z�|�����{J
r09��h����A�982dC�q4�J,���?��Ց亩����Jy"])�%�WV�G%E���>��,'�!���	+��A�O5�%z���}�l��Ɔ:�9sڞ��̭��\yg}ENN�'����
��fq���@TŀT�)Sr[}3���v�DM;���!���D��Q�W�@ebC��X���F ���<7�>���2	 �&8֡��b�|Nn�Rb��� �����2��p`�S�q�r|�_@V��s�1	�y>�'_���ƚM7���"3M�L���3㣬���l�t	,d�S�B��x�+:�����)(�e���l��c��.w�_�G9q%�x�\$x3A�:���#��~�=�&����wF��E��L�)��KŠ *A�Z�#�F�ɣ� D�W�h)Rs
��CWR=��ik@��"|��~�7��S�¥K�%�c�r��5R�v�]�>�}Y7:k�#�����
$�ʬZF��y�|>�z����n�
�  ��(`�u�꺵k�3���`O�>�6s�����\���l�,��0i����0���׀��(fG�3
�cS8u��C>�S2L|���A.$8��	�L�e���8���h���><Ĵ �*��b-r���P��4�S��s��:^��w,ښk-_��w܂D�5�*��D��wD]}��VW\,��s��>=��4	ə�/�@ɼܗ�}�H��GVN1ҳ��h�����,�y<2�qӦ��Wjm�4�'O�&(Ϡ�b����"/;#=ظvV-��A��c'p���n�r$����R�&;tI'�����"��n��%c`�h�m�����b�E L�<��Ȟ=n�- 儠E��F��O @ m��A��0F|K���э��^tw���w}���Ɛ�p���Gp������� d������5��hk�Bo� _;Q[W���.���hoo7ӱ��^N,��m����zѬ
g�̕�_�N$~��)y4���]��m�E���-2��-�H)����iCcdP#�y	��)���G��F���C���E�Q�L�T�)�#�K�$O$���"i�:^�<<d&<���Id����|7����1�T2L�,Z^E�G��kx��}X��(�\7�r���N�2�0�)-+˒���dC�)�j�~��36�{�=�]H�������7=hV'����U��܈%+���d�l���݉������{�1���!����^:^���}3�uD��Q�|[Lɉ0F��$��T�dM0R��ƑI��)8IrJ:���u�sb
 73�}���#7����(��lf�H-��X
����U�g��q�L�,4�5�D�IOVJ#���� 'H�WN&����:F+�R������S��ზX-V�|&N͕�r���|�	a�?myyyX�d	23������ ���i��p�����i��!?b�!$��S�PU���*p��ضn%nZ���ǲ��X8� ��(�HB�;�ӊ�?J;J�F�47�6�ΰT㎮�C~���n�}���X��!�.�����D��#���;�#������)����Bc�^�>� �0LQ>H�V��Z�(>hC]��
�	�^���	����s7ғS��^x�%	�+5EȌ�5��U�����c$�k�oDog?�;?����\��f8�(���&�����=>o���D�����a\�m��=���~�r��u�P�dz���n~�Fm}j��q�r+.\j���8w�-m|�y2�DLN��lg�&�����HqX����F`����i�$�/((Ek{��)���s`�%(>��z��Ε7J��D�4
��u�u�����$��Y �J�I��"fzɮ(g�beE)6-��*�Vd�"�E��`�;��p Y���I�C�;
�I.�g$#+5	Ąh�ٙ�ၢ,Q7a�� �oT�y[�����A����#���&=-�2$���s��Fj��	S!����#k&�*oRB<��1�5�斕���n\�X�n��j���l�~�͸��p��-x�q�M[P��k���ޖ�)�l�U� �qE�OIK�Ulg� �X-���6^E:^��(mf�����6��P\q	M(�BSr��[���y�ͯ �.EFv	2���;lN�,Bzf�mY�x��J�Q���x����c�P�fh2��d畠��

����'��T�7ɩ��id��d��d��f���?`Q����4�����\��ŐL��E��Tz�kQf��)Z
k~F����SݣQV���%X\V�B��Qc��hF_k�:�1�B�;�d��9i(&Ȗ椣�(��Mq^�����4�4����s2;-P�@46c��5�9���"Q�\1Q�ߌ�c�1�ۂ��z�[1�߄���]����Nx�n'�
�=���(D���S�������a��Ԁ /����[o�������nCA�ۢ��l�ZTV-f�TDde�ݺ�ׯATЇ�x�/&`[�GZ\,R)�)�'����+K
P��J ��x�,��V��X���y��CSd�1��qV}2�s@<mYe4���v�\RFQyq����������EЋ��?A�<� �Z=<���3�)���lX���&108���ӛ�敎X*Y(h4>!ޞO$��\�+׿H�vV��ReE��~��J=aV���u���ID|�2�0�<;n2@_7�z:l�)��o�ǅ��d�f�#=�C�����[@����\"ɶ�>����G�&P�0r��G���%�����[m���Hy�#���a��-�_� I�dk��P7Yd&Ƽ��ct���>��%}C�:2Љсn���C�&��&��t��E� �#i$-]J������n�`��ؽs֯ۀ�5u��K�ѓ�����p��q�����܈���tc���^�C�z�k�u񓭎bd��]�{�n��1�R*
�{l4���Ó(E�R�{i�&�]�b4Eo�	� �*m
�Z��65�UK��+�:�D�+�t+ʍ��)J��k����.�I��8�eff�����)x��AnN���J7���� �������K���������(W����d�/ףdq��DJ�3Q����#�	�(�1Y�3ғɞȲ����>8�F�#��]��QĤQ��"��p�p�s�j#6z���5�b��r�s�vē�8�M���v�:���6,Y���p�"��%�����W.�F���f�R,^X�ϥ(*̶��W�0?iI($@�+-�HS�d��ɟ �0����#��Ʀ��ևw�ų��@SS�U�Ǣ�K���M��8�C�"LƝ���X�za�#����2��eZ�릲]=�Q��+��[y�Q2v�3�-�Z�Fi��aC��I
lͲb~a��V�d�}��jbrfb������:�g�z�m}����i1I3���+�^%
�b�X&��z�I�T��E�Ѓ��Z��������ڜ�t��1�H�a$�)%���X�A��#��i���?}�[����yXVA��Dc��cã�MK�L��}����S|K��d6�ar��8��e!81�ξ!�0�J�}�N]@RZ�c�17LOEØq$��qpϳx�����_�R4����p`� ��̗�Y�=�=��c����6��(/�99�w�G�-E�q٭�yIUb.�T����}b~�m�xv�Q�=r	�Qeǽ(,�GA��F_� �k�@�D����mX�i)r��<҉a2ͥKV����"M)�����L0U�7!^.��>�}��d��s�;8���y\��6Hă�`�3�r:*��ĕi�P��ɓ��TE�h�elZ���dL���H��{m�J03�DE돥Ġ4��y� �Ns�AWg+r�S����,�u`�nx�#~�����s�̕�Y$YɳP@1ĿV@z%�$/6�ԅZ�RO!X��e /̓I� B#��LKCIa�EM�LMs�q��6a�E�Y��`�L22�xn�
�Ȗ���&}��d-%�F�LԦ��f��R��*p��m��4�$F�Sx�buGG�K����Hv��G���h(����
���q�d�.-����q���x⑖�AvV.�̏��Γ�NZ���:���Q����?@�`��I~�'NÙ3'�o�.9r۶m�����H9�ŗ��r�AaQ&�2-(rjZ*�KB�/.�B���W䣔�]^9�uJ5{� AI6����Wj�J�d[+���-G`�g�!T4{� U��_�+&���G�K�@��We;��$�GA)��S���/�T��p�{��c��~�n<ĉ��}������c�Mb��j��t�\�"5��C�}Jo���m�E��-���sL�h�!�&(}�EcQ]U���l�(
z����=��%%��Ka�t�f�A��*JKL�O!�)��%�Ҁ�57R���K k0�6J#U�x����u#}#�HOIB~n��%-�������O��	ngΞ��S�p��i{=v�8��8��g.�RM.�6�܅F�:s��/chxa�'��Y�h)���B�]y�`V����a�H�jV&�rr��Wh�Zl���6�и��C#Cd��<��ڋ������Td��5ǕS��Mp\�b1�ҒȖ)&c�̪�	PP�?ٳ��>��� �A�U��������$�|&a�U��}lK���{ȬK��MI�_Q�cx��$'ʶW��^P��(��(�<�]Ǳ�+�c����.3���&��=H� 	 ��\����J�g��,��5*������k�h��'-a�¥˱}�2��&�t��U�Y�==�BZĐ�QN��	x���DX�+C����x�s�!���;�; �h�_Ag��Ғb�������n�W��9[��!�t��>�C�I�lZ�d)��݁�܀?��� ?�w <���ݳ�uu�b�`5���599����u���F��?
��Qky�$x�����
��� �:[k����z8a��m�� E�֢��?+��D]�����d��l�QD��t^#��� Yd�����?���N2[�'���.����ѐ_�fT���I̿]O��2�v"R���e���"�ة��ɏL����褸�ʧ���@_��S��1!�K��n��?}���Ɲwn�I���g+���͕�r��(�Ҋ+��ҥKMGz�
E�OF�����:����+�ˑH�4��f�3ٹ�hi���ٹH�x�Uy�J� wـTZaAN� %}�[�pg7��~�S��x��`�`�G�HK�@@RDv-6-Z0w�~�QQ��r�z����⸇u҂�捫)nǣ��?�ɣ�t�1W�Ϗ`@lL,�f(��ʲ3%ƒM����-M-��f�'l�	��ej<�p���O���~c�>d���=XT]�7m@a~Y�q<���xꩧ������!���8�?���F���x��q������[�W���v�؅�v	%��Exr��gy���
�|���<��R�N�$�eѲr�Ґ����g��I5=fvV��e�}f���S݃c�|�v/���O,7�]Oi��5������[#�#{wǻp�=w�����2ԏIb�̕�[l՞�zjJ*%�B��k�U!#��G4.���[?z-m�X�~#�u=��#8���f`����oj�XBVv�%`�
�͸ܘd�)��js������Kː����{���p%��?}�I�)�O�X����3c&�不����7����1ב
� >�{GSK;���q��I��=o�{����H�O=�w��k�R�\�nWp��%���S��*3+��x�y	DO?�3��x�v��0��h6IV�{� �ӓde2I"�R�����sH)��~�X�w|p��Y|�����PYU�լKEe��;��D��0�׏��œO<A�;%�����;l�~������g�{�\@W�^�͛7����:1����(..2�%ٓi�|�4Z���ɔ��r���%|�0�(�L���-O���(��jEL4�PvW�f�x�%�<��"���R9{��E�*.�ǃ����Xk0Fߜ��y�\se�\�"�Y�~X�b���ת\�Hg��3��gk$P�+����H��/���I�ʞ�T����X\n2��8g������u�@��g��ƣ��	Z<�DGW/��s������dD2Cjm���d�w��HEpD.e���lu�;:��o܄���,�������s�(.�g�Y�)��f]�LOCyi	�23��`��VG[��&Њ����*�硪b�銧'��s�M��QZ�C��KQ�ӓ2sJ��k9	$��a����/�WTc��M%�	B.~7cls��0��-h�i �ss2r��{�5k���U����J��=��}��E���3>ߐ�Ĕ�˽��ݎ���ü�����'�q� ��NNZl���%f�xa5֮Y�ի�cٲ�X���%E����ē�d�_���l;�7)�^�5��8���`���P�Y^U�����{Kl�̕�^;҈�ȁ���^Uׯ��)����9���j��\�O��iRE�1��nEB'0X%��4E����gZ}�"�6��QԮ��G���|���#����=�t�ZqvD�֖z����@*F��0�/�އQ2;�}�����-�2XN�>�zvZ�о�8��J	�b/��ቀappJ�!fv뭷�mo�	(�o�;��<p߽X�x
�q�捸y�MX�</��8t� A�[o�	�6n�l�5de-�ͼ��3����R�Boj._��%�8+�a߾#�x��ueq�}�����2
{��,��6o�}�ߏܼ��X�N���l����^�<A�"N�<�s�Þ=����><pǎ����q��	�:q�^�Z[	���C_�N��c�X###�6q���т;756Z���Z�tw������DżyX�j<d��1�pܯ4ٮ�x�a͕��(2�Yˢ$��%��^�M�@J���^�LR���Ԅ^^��#��Nr#���#�X�����!�4:�L���(��iٓ��1���8��	{����E�FjZ����:n�#�N��S��Rc�@���61S1ܱ���L�Nc��
b��҄��/b4�EZV�rs�D R@�8����X��z	�)H%K���8�̠zQ56n��m��$�(?�<��;�p�֒�ݸ�F�r��"�,[����hnkE����܅Sx�ŧ��Ǳz�B�/_:�I�	��A���[2>����4�wJ�ȉG�����(~?m�aM&����9����K9�	��ed�9y����\kYd>�
KPHV��[�̌lN�N4*ٳJQ��ޞtut@y���V,��d�~�Y{il/�j�v��jt������"q�%$���:�\�+o�"�q��DB��dVe� �,���ʕT#���~/�^�G��ԝL�IKDR
�ED�� �A�&&�^����qG��Nq0)����@���-L�� L���FcK'Y��Ӳ(�S��KH���x����:,&3��m�6.��ґ���.(����pӍ�`~7mo)Ap͚�f�S1��2�����I��!h������ˇt�����b�ڵ����K���6}��[��9|����V�W��)O�c��#�Q�B&�n�z�����E���b����,�|N ��܌B��^ܹ�?d�]v�-�PZV�	f�X�Qn�� �������;e"]�tV�^�{]���U�_��׮�M�n���n�m�߁����v'��|+��p6o��7g\Ϝ=�̬l��)ެ�T,2aK��"�Y�y��c��uذq3�s-Z�<N��9d�d�m�뤵s�z�����ru��;�\�+����&���鵈Azu�B�E�P��Eh�5���@n��Fźv1�!�&�I��$	7ӟ�-��Lpi�>D�8�1��FGw/�Z�n��qB�q���H,U�MF�DA��E�܂bL�G;�}z�A=B}>�%�4^���g0b):˿V2R�	���$ϡ��d -��@-J�S|n!�T�Д�b���p�sV�*#F��)LNM�猬4N:�6�UW/����-꼊��^i@���xm9H�e�L��B�u'j�x���q�C�y���{/=���, d��ݪLl��m>N�"u�'�Xh��	�����{]=���F߀�^Ϝ���N�k}c��Z�B�|�A��KPT@���(8R:�+�U���0�|�Nh;P����D_�\����;�s�R�c���]�2����ۉ������EȔ���8��\,�����0�����G<Na^u:k� ��Eg剿��b�?���Q�� Y��]������I!��`�s�����QH����]O�M܎o|�/!�%va���0��O���������G��1�g+�����Oæ�7������ୋ,"�x#6�� :	R2�?{���oc-��?�!x}��N�8{)eG��ބ��|�>�>�O`��E���w>�;�����?�q��}�`2ݦ���l�F�	Z��y�� ��g�y�Wwq_�����A\�x��7�����W��_����?���=�RR9q( 3�� ����yP�I2f9H?-��|c����>n�e����b�9޳��4�XD���hyϜyn�Yή��b�`/�N��K����~7�c�鄏=DQlVO��Z��\���C��}���^�`�W�+���k��3�0�;5�L'���q�h��r�)��ϏAE0"��A���MN�aN9��ɌF}A���j)�G�q����̦b�=�OH��4�[%8^����(�+��������:NL���3����טPY���U�O)����Y�Y�a[X!w$3M30�l!������������(�W����@� @$d�#�u��'�z� yݺudf�xꙧ,��D�M�7�޶����>ژh�����T.��2闥��H��1)a�q��()+�y��܋/PtnGIy.�}C�����ꚰo�A��w��ǉ�g(��A�?|�$Ξ�AMM3.�^�܀���	�ʤ�ĭ�>��Vpҋ�('���!c�:z��Ԇ��v46��������9���uhni�=����p���7mڄ��T��5����$��+s��	�Z`֊���C)�(�
@d��jnB3����\}j9��IE���\�q����w�]��F����]��	�$�&�Ao��F(�������Tc�ZXQK�Ɋ6$�c��뫋�/��4b�a��BX����Nv�S|_\\b��C��}JVߥ���O@�EOb��OI��R��Ԫ�����;�˖/g}��#bt
-�^C��Z=�r;H&^_߈����_d��i�f<������0;Ny��U���C@o�XG��غ�����j)��d喢�j��؈Uko��P�`�/X�e+7`���f�X�v�߂�7���+�c�u(����6�L7ťըZ�ՋV��PV��γd�z�Z��7nō[o�֛oǖo��-7c݆����W�<|p�ê	&ȉD*�*Q;Ε��F("Rʞ+�۵.� .� I�EwWT�i��b���$�Z�p���$�	�xPȁ=o�*U-AVQ�2󐐒Wb2��<��M�9\�'`t��^��l��%�L�����@����S�e�ƫ�T�N �Ud�O*-�b4��M�;�j�_�J��Rgfe�<Q���$kBPa�d(������,���Aܼ��
��R*wX9�DF��(R{|�
x�E%�� ����&�Ĥ8��tã##�~�D_r&E�w-G��@��(0��	���\�i����H9�\�:���r�!ƕ���X~?p�F6����W�� ��0�-}��3^��	�(t��o���)���B�a�#��K<N�(ݫ��x��@U�f�̕7B1�x�M�H����*Z������r����iW"zGB8p���w�Ԣ�?�O6R
�#�l)*>	py��Q�ډ#���ȉ��Tۀ��2�����'��h���%����+���L����W���a�|̵��L��s�fR�W(�S��P��5�'�#���VjZ�5��9z������_�>���ⓟ�����M<��ؽ� ~��������O�Ӽ����2��$<�Ddgf����دTy1_�_�ɕ������-���*-��4�g��|�����$%e�}\l�&L�q)��<�X��ڍ7;�̤q���9@0T��1��t��"�h�a;齬'��?0N?n���O�blZ���8�XvQYJ�����ݽ�[144��Je�V���9jAp�̕�]�#��?�t�׸�A�V�b�m}8q�a�L\"�b(F��s)��剖�gkh�@mC.74���u���khBKG���7�w��o��F����IL�}���@�E���
{T�Dۚj�a�Jlۺ�t��:v1�'�|A��V��]�v�r���&~PRRveq������=�D�D��S,7���c��p��Y�<��P����M��/�`��C᳸p��v�����K/�ƹsLu���c� ��3#������ϛ8������Z�ߗ�άoG&e���ػw�9�=KGZTTH�
c��c�Q6S<�i����{Nf(E��J�t�zfj?yk���g̻�e���#��}���[�XT��L��!'~)�)c��I��Y	�������K�|�b�{�������{1=��t͹2W�u1ҥ7��{�ob��[���Dq���k�'g=��kO��׋3��1�F�;Sd��pX�#Vp���F(���������?8B� ��w�R�Fb)
��U�P�G$���lv����X�b	�ݴ���:��4�}~'Y�223-h�*�tQ��1ر�%�͗�=��3���`�3u�0�-m�T�������5k�b���f��f��n޲��~n�~n�q��v��^l�r��Ya��j��YC�X��5�A����̂,����;++�ǀ ��+O����d�.|���<���Qx��]� 5-��N��$	�rkU���+�����l2R;��F���;����0�^�H�f��x��h�7z�M�Tb�y����U���W2�8s#mkm��Eո��v���v=Z�UY�m;�\�+�b=mP��#
HE
8.��(ʽ����ph h��x��Ř��+}�+1�9��.�B~�"T.FA��V ��)�yH��Frz<�N�'Y� �aGc����k���u��Z��}<����Ż��t�:�>K|���={��5�7����ᮻ�F9Yc]]=��A�)c�����`p�]抹z�F�W#��������m���7���ތ{|x�;p��{�~��(�q����n���d�!8�$��&&jKA:�0))��#d�uy/E_������I�$wccӣ�:lQ���ޭ3���ң8�(Ȳґ�iAks�XNVQac������[�L�����|�����T)Z�R�~��U/P�g���u(�F�*s&�r�m;�o���kM��rYMF�*��"G���;]z�̕�_�A�(W��H���CFz�����_��V��b+<@:����r��"��ᗲ�$��<��96\���1�􆺎N�YClS�!F���QX-�$#]�r	n�a�cN�_���v�&Ql�EG[3��c��HIr#--�w���?�C���/��cǎ�j�$̙J���L���܂��P׌�F�z�IW����=�q���;p�̏𵣫�̱�.ך*�ȑ���Mf����g&Q�y?}�����3��2�ںZR��&��﮻�@qIu�=��Tr&P�~�g�Vq0MFM��%�����Dl13�g�cd/Ʃ�,�;���ez��z4��R��${�~6�~j*�5�W��4śu)Z>�$����T����ތ��z�$��哯z:ϖ���y�̕kY��p��W2R�p��J�w�˕0z������c��NFLZ&�`�Q�Uy2	qs��f��(�����@���SqP�8�V��C������h�c�
<���O���0���A<X%�]�3�Ї��}X�|9�|	�߽���FA�C����_��	��GW"X꺺K�!k������)P�,+�)�FFQ�F���?]~��ϜE���cز�Jm-�d�'���df
�|��y�"�Q�}��Kv�	���ҥ��/���yi/��K�������4�O��_�倢��SL&Q	DM��S�!vgb3�\�5Ϫ��Ԯ�0���3Y�%L�֝�K�MfW��x0d���)�L����q��@R�\s�3L���ҋX�����DuU.\<k�T]��v�$:W�ʵ-�^��}�y�>NL�z�<s�
�t��kn��BF:k��A��+��fL���PT�!��y���{1U��`ŧd���i|���qf���`U5�z��=��@W�&��{7�U��m�X�|1nܲ�m*�}CL����"�FAa!�:ZPVZ��V#U���2;�Ea͚��:��ثW���U��q�F,_��
�jv��]gp:ɹŘ�q!8��e�u%���U�WQ�q�H���c~�b�܉��|���T�nŲe���g(�'���9�����+�̍U����5kV��މ��4��;	�cHNVjMH��?����hi����&��������|�A�8d*7�g������Q~��F)���<����;�t%#��&q��wݝ���֏����1�ߎZ��ё!�)�Jm;�cM�WM�Y�\�+׾D��y�JF*5�bG����M�2
�u�?{����&5��t�B�Ź��
9~�S���P)FBҠ�s�^b?Et�5Kx'S�:MW�+]!�i������8(c�ǰ�Sx�[�������9�-���������"�a�F=��ް����� �nF���)a��pcY?����$6�l�a�s�vE��Okk+~��^�t�,2	�br������������hklZ��.&H1-�Ɏ��������%Y�S���A����X�҆h�]_b�2}���BAA�
r�Q����>�12��Ti����@ �yYX�|	�[6 �)#���COO/�?K+�rJ��X�R��a������7^2���~;FV2˒��X���t��pPn,���wR���^(G��߇���l��ǥ����Y�+=KeG�d:W�ʵ.�� u޿��*�����]�r�מ��.tQ�߁�Y �`�0Ygx2@�V��$fdv�I21��S�G�;:���#�N�|�yFސ�Q"�~�$w��j��#RiQN&b��ҧ��G���>��5 e��}�3��?�8j�[-�ѡ�;�y�
|�FiQ�.e��O���bb=wJ=�WMB�˛�F����ѳ��N�)�����ݳ�s�FP�$������>20�h*gkC=F������[M��5�FV�J<��Y�߫N�'��h�'gO��#�(�0in��v�u�vTV��q'�����^�����1��}kdtĮi�Oɀ����ZĒ~���555&�WWWY�p�r�BZ�hYb���x֏	V����������P\TH��X_(���C144��2o���\���i&Ǯ�T��׺����t�}�K@��8A֕�́G7D�+�&�ab�X�U�i2Q��b�V��/J8A�F�i�I�&�z���hF�J�'��D`j�â�J�^��8-`���Dc����;�h|ђ��`�˗/��Mܰj�HAH� ��*d�$������q��EԐ�z�d�D0��*��
tuw��PRQ���b�^�
7�Ö��|�b$��*gӪ��gO��.�ϳE�R[�:��:��`��=��³��. ���׸��;�l�BD�}��/�������x�3�ONN��K�1���f:��82��1�OKW���|ܲm+֬Y���N���LCFZ��R�X)���=?A�O&:�׋SǏ���+W,��=�v������L��g�E<��lcϕ�r�0$���^�AJ�E�d�$��Z��c�C�ù�a|���=�;�� :��0"�)*���R�W0M�	���fJ3a"�L�P��I��H5[�R���f���^c.��7�"knz���4�����>�~K�&+R%���Ù3��r�-�,v鲅e�,/@��X���t~�5�s9�m&s��N2ѓL&淕��wB���ժ�eE��dub�Z]׳���R�<�(.F%<��_3^~v&��V2o1x�e9�\��<��S��C���4�s_��@X5��G���`��q����-o}�s2��ܿ=]]�snC8w��2����Hmm�EMm3'�!$�$�ZC��LEW�+�\ٵ~�>d[rR�u���q+����0������U���777�q���_��_s"[�(2]=Ӧ���yc�ڤ���gM?W�ʵ.������c5B<##͠t�l��ߌhϊ�h�v���}�E��wF���u�`@U�Q�N4幣�K7:=��`�)����(��j�^�ÀT�J��dl����� i2YY&A`�g�w�L MJ�s0���c��O��kڰb�:�Y.���^@��o��u+vm*Ϋ�yZ���KG��DO�ʇ)O&��EJzAB1YY/��y>�t*�\�Y�ߏ���!e��7$��~��!��L�^R��'���IWI&* ��C�XR�G0~9>�g�*2�xwE�Q<���p��i�^�����#�y�*�/@<g��nE��"�QEe)g�s:��@EE�-�)F� 1/7����*���
|�8��;|�(�ZZ��D"o,�}^�x}������O�����Y���ԌS��P����f����\�����T���T�F�u1 UU��wߥ&��L�H�8�I��v�q�����4��C��̠de��g$�#%��'�@V�|���G�D�8�����w߃���,����͑�����~��X�b����nk��#���q$�����̄��vM�:۔ٱ���Z������/%Cz�"T��Xh�, �@s�/��l|�?�AQ�T�c����P�F��^_���DL���♣�&ІxOZ��6�&���D��
j=�6�s�7��8�ʴ��|;>�'!X�Y��Za�;��؄��T3��sE!7;�ť���EEO#6��=; >Cv�D��UA{{���mذ�R��|Jn��f%���	���&�;*���8�p��A����gYXsn@C]���҂�X�Xid�k�̕k]�z� � NQ�_<}	�{�%c�O�^@:����,���e�(�46�,�Ӏs)�OlT�O�h��e,���Ӷ�������������#��?xA���b�g.w�O>�dF>�X���M�b�V,����Kɖ2�,�H�, U`E&R�:�Q�|yA�]���D|�ʭ 'kzp�i�\Z�SS�� �:����k�F\��$h���	V�Q̌����:=�ŝ�m�+z6W<���j :J�g�晠��I/�6��O�2�[�ۮ={̴��� ��z+�2���;q��Y,Z���l�I��>x�x\3��B�"0Y��O1�|��ǲ�����Ʈ]�,VA27UPm��@Y$��!'7�&$-h�QR(�υ�7����1,^� 7ܰ�������55橥	�YhRW�+s�ڗ�Ҍ,�oh�ހ�u� �=u�~����Yp���D�Q�+�����NX:m3�i�x��bf��d�X�@�	�!��N��������D2�������)����-�r����V|�S���D�����O`��*|�O>��K9���?65�Nbesn������!b^�Ĭ�^���ķ�R3��h���hO
���db��w���&S�ARB<�GV܊�����o�[ڎXi�<�4����.3R;��1�=��V;��
H�������?~�"dmش��Z�Zٍ6aQu.��q��p�K/�֙J#)1�,�e�4N�_jZ��}	���S�Tm�m~�MȮ�$#8���QA@/s1�����8s��~��n�le%[ҋγ�L���Q���\�������l[����Z3���\��҉�m��#&Ai.$*Kǧ�o
���&���'��{��sL��.4�f��ݬ M�b�
�!���Zܱ�f�^�����̈́֎�ܹ�����s�q㖍ؾm�S�&��E9Q��U$�ސ�9k�+�(�x⠽��Rm3N���cy��d�!�P��s�>R~���<G8��w��ݧ&�1F�&_����A,Z��dO%��"%�nT�S��xn�x��q�	MJr�<N
gN�0��w`�X�:>���!��T�wƳ�����GQSӀ޾ax�Az-`LgW�[���?���n��p"����a�K�!9-��ʷ��4�&�Ѻ�=H��W���!3 1)��3)ז�,Z	�'N���[�l���Jtp"QΫ�申͕��+���z&�PRǜ�<�l���* .�t�bS;b����B6CP�~-�((��Q"��>���G���Y��1 �g��a����Cg���Dt���Ȃ�'�?�y�6�Z��Ω���3���McC�y?-YX�$��X ����:}gΜ2�S:���V��֚H�ܳ���C�q������^��ĩs�$�cY'eE���O<�&��.`��·D N ��G��݁��4����L8Nq_�A��R�(��*�K(8IZ�4EH�w�BPÁ)�=t)9�\��OǍ�h7�4�@���}���8K� f��8)x/�ER*�S3�}n�bR:�T2U%��dEf���f^ZZ �~wB�Y(���J_��3Z�+�L_����P�����n��yU���=�9�\�͖_��	�9���Uq�8�ǹ�h�)<��\�E�IH'�
<s�lq��Q.y�>�`-(M�c�w�Pt"UU�щ������w<V�J��0?$���dk�E���c	ғ~�z�g��g?�}�9|	��K�A�@����z�R�?rp���o����f��������x����(]uQM٭�QՠU�,��������q�%֘�W����uԢ��BA��2�)��;)�L�">������I]�(),�≈�
���������+�]����|o�_[TYL,\���4����7?���4�������)^�@���9�z��9@�������,��0�-J��L�5Y�;�Q��Qr����D�Lx�ׄh�C|.�]��C:d�D.e�$�>9Y��O�4��8}�(֭Y����_"�m�g�N>{�6�r�+s�7R��"����']}br
d"XZZ:���c�nZg��ҏڶnD��@9�'��,�X>�Q��L򍟚 ������d�O�^�bbr�L���!A��&�"�J=�"ٟ��e�Fs�e�|�&�_�R���b�~��g��N���c�YXUn��;��6Y[���q�%!#3��23ұq�F<��C��N8��9X�l�=M�kf=��>���s�!�����/;'�Dw��9������"5)�W��8����r�m����}��v�blZ5��Q:R/���se���ւ"/]�y�EN����C���I�`��L�N��*ށ>��,]:Q���N��5��zB�&�Vb�aD�%mH�Ф$�M��b�3|���q��ÉE�^��0E��*'��X�̪�%"���d�7߼��<{��;)1�~c3�\�+���*��y"������tbƵ.��DI�l��և��6Lǒ��%�T4 �$&#y�a�?�q�gx�,���F,v��e0C`��³)��,X�\7ȋ��p���
P�X�������l݂�d< �t��;J }I)Jk!�� �l\���"��������r<�ЃX�z5�)U��X�h��k� ��R釕*Y:>�C����0d�d^$Q�;2@��ţޞv:��݆��N�(�?|�=شn5�"��k׮Aqa������|�{]�l9���X��RU���%W�͛7���~6ߋ�`d�o"�@0���"~O�'9��y�ɤ)<���
#�N�@�1q�+e���,�5�K�V,�âCie�lU�q�҃k��	@��5fd�!9)���z�M7�X���"מ+s�P�����n����ʮE��"*Ym{?.44c:*�n)�	�@t*H1�H��AFj"��1��y~Y	�g��ś�|�|�	��')K6�$�0Y�S"%G��F^,��5F:e�F�fd���Pn�
H�|�9�'��ZӸq�z���L7
��I����i�=�l0�4+3Ә��)ز4)�Ҥh�gN�Au�<����[��0n�u6mX��Vុo��w�N>��dQ5R�d�x�{ލ�+,�IsS#r�s�MƖB��!�HO30ҒYrJ��b�������{� �d�G�֯����=M�R��<N"��Wg��K�D�6ZY��J}\�T'��p���活��*6�	��O�أ>K�WK[<>3%�@+r�&S��J�(,P<�V���"1�Ͷ�0@����ε��\��E�Ҍȑ$26�U1��54�<��'� �de�d�3��X,�(�k��ͫq�M�p��q��jlXV��.Ö5K�~�B,_X���\�x\���Ef��kQI�Tn�6�8�''w�b��|�h�G����"V ��V��Z��~�՗�>T��������M��;/&&WI����Q���oن��k�*�W�7vi����|3��ַ�C��{������r�����I�]n���l���� Ã�d�ݸp�^x�?~��S�ϓK@���<��t\<��@�'�,0�-04���1x�R�Gb�7��m\�\1an���̢(�},7���FIA��Jj��8�҆p����EG)���曒,���-�)
�̴, �f�(O)�C�I(.&��(�(�ȖC������8�8F�u�^o��k�tX$�8d�vFS���J��b~QV-(ǲ�B�&�`�ߏ����0>ԅ���S�OO�<[U^���\d����|a��3yE�c���H�M�,v����b���C�/3#!��,5##�y���iӦ�����o�Sy��X����Ou���ƥK����-fh�ԓ�O��_�2�q��XVg{;<�T��c^Y�s���Lv�v�ux!��Z\���@d0��A4�7X�|�p��{	HZ��5U��x��@x"��p�2�'��c�k���z�N#��=E�H��# ���3�AD�z�S�������Հ5�k8���i���Ӽ�d�!�N���X���n)���e?
����y*5�b�
D�ƈL�se�\�" U���
�"��9%�+�P��Kpl�d�`)�ޥ�K��B �a������Vw��-�r��� K� LM�CNf

r3͕Qv���?.�W�hJ"��]fFW@ƫ>�l��~�t���*��@Q�-}�2{VWU��������3d��e������#�ҊL��1U����X���׏��VW��!86�&NK���KX;��(e��$"�ׯ�������;�4��ҏ457����Jn��)�+������#�!ۜA2��'��m�$��S/~�@T[��v	�����s�z�3��)n
>�*�O�-����*�����k"�g;��{a=����6�q����.�zy/m8v����mfh
��	X�[�j�̕�_��k�*W�r����V�e�>>FP�Aya�U�#/-��n�h��3�P����T7�S�G���J#� -)���(��DQ~6��C�� �j�_��ɴJlR��jJ󧿯^�U[( �CW��9�|�NU�?��O�S�$қj`��.S�I���S������� k��Z��_����X�zOc6���#4	Wy�d��������s��P��S�w���X�d)�Ȏ.\HЏ��-2���8�2�R�|�e�E�^тU`t�7BAt�@��T�����:�������@��=fQ��7K���v�ubd���8��G>��Ntw4�������I�eY�D{q���isvV�1�~�WjYGtD
r�UԂQw�c`���� �Z�\�+ף�I�]�5���6��}��T#ܩ���Ӱ�*�L4�|]mMf��E��.W�Bt,��o��Kv�[T��B�2��l�;�GbB2*�:EV�hv��n���7�^��wކի�d*��4����ݎy�L��6oؼ��h,E�aL�i*�qwo��H*�� Y��_u|�5oD����@6�� ΟG]}-֯_�eK����qǋ/�����)	�{�z'�+V:/7��-8u�8n��f$�ቱ5�4"�(Ϣ�[�x������p��9��8ۀ̜u��m��c��e��u�Ks<B�=|� ��.cx���0�R��p��v�QT��e�`�*,\TI�����l[�t�E�_�`>A�K�, ����e�l_iI���<G#//����~��K�V.�[�a��%l�l����o{�J��#/+��؃��[o��z�8YLp��VF���o��Ε��B�fD6�wy7���Z���٤�Y���������F	�育L�d�#�ߍ��l����L,A��!sA��e�42c�*�����M���e�>J�F�˃��B��\����5����x@��9�5$��d��?���)Cs /'�2����|C�V�_����)��V����������j읻v�-�m[Q]Qa^P;v�H�>�e+�#3+�`�D>��������k�����a�#� �)�f�)�uٱ�)ĶR�����M�q��E[���]Ѹy��5*��C��O� ?=ty�=�v�&v�_�lY��7o�\U�W/�n�֮���k���V-�ڵ+����5+�ukWپ��hn޴�߭����ha�rYf
(A�f��`au�߶� �N��X��%E���!��b��;Av���϶uaR�,s�t�\���7�ɱF�ъn&��kYL�Wd)J��]d�)]_vf���-M�H&�(:��9�&��P9�$f'y-@p<�X� �=b,�+�@��m��).�-* �#��^89@q_���j�sF�H�;m:�)��A�Z��9Sll���8q���H�C�=K=)G��Fދ�ad6m�2���ee�7��n"[�7ଚ_�B����K����̣2���h>19��D� US�?e��\�V���w�E��dn�d�J��	)���� X�IAV-��,���#���۰n�l�v+敕#��Q�������PLoEcC=j/_Bm�%�PWSCf[���F��Aw������&��d�[6o�Ѓ2���E2�'�|?y�Q��{���oij��ﷅ���n��;nü�r�[�1�U�̱�$�S����4�Ε��F(�p�`�m��H����f\�i$(x(:V��0��ntvcIU��+�zOo�1�d���T�� e��,FV\Rf~ݭ��E�wS���u�8�&�L�1q���޻o3��1�r��w��^"p	'	6��uۍ|� ��O~�

��a�Fc��ݽ�3�!pcbm�"��pB7�^�9�{E2�z89������Vᕻ��F#�I��7nF!z�W(�ޫg{G���K�#���ζ %�ϴ{�^�/�0��wl焓���<��3d�c��m����cUݷw/^ڹ;^xG����{w��9w����8|��>�cG��8�;y�$Ν=�ӧN���M>7l���ё457�����'o���VK��|��6�,^��d��l#���#�AbR"F�#���rqIM1W���(���ˎT�����]� _@"j�>߀چdd�aAu%J�3��Bxl��#Ф��b���'1I��r�8�O�:.�*UU�.�B��Q�ťU���m]���#��&9X��J�	2�e�g���f�l�W i[� �{~'���-ݨ��2�)�Q\���6�r~��@F�;yY��;�����E3ҹ�ȺNd�R�Ο#Ɓ��k�.�۷��>x��j�K/�m�L�R�����m������t���M� ��2������3Ʃ�x�p`�A3��% I�q�m�"7'��=���|ڢ)�Q|^�h�I��FMu��x	�KZ'�Bdef����1�[da���Z����)tFF�-rUUU۫�$�(���v�QA��d�rNt��9	)@̼�J$��#j�'�-�t�N�GwO���uV쥧�Թr�����X��_K�Y ��O����ҍ̬T�+EqN*B�}�������H/Y��<������Yi�Ri���\ǂ!�@�R��ՃK5�&�NSV�xe����8@����:�}׭X~He]I �ĳ�퀛�-���)��둗�FF5�s.S���P!�ɍS��`��{^^�1BE\
(����+5��I"�V����D��4���U$���߬d6%p��ĺ��q�mwX� �����iO����61>E�l�bI�q�h<��nc�:�� �r�V���`<8a*���G�D��e{i2H'�-Y��Ȅ�m�7ݸ�o��M�q�M�p�M7c�����ƍ���K��n��\�%�%���g�\U��i樐��d��J�[F����' ����K1ĶQ���q��)�����9wt�6�����K0z�:�\�+�r!>)Q
�ȵ�n�u%� ;<{��]�HKKQ����w ]-m�!��@SIN%0p��BZ\�%8(+MP���������NL!�����SQ.c��.7�	hZ�R�(y��v�������Ү�<���d�Gx2H!8�R���Η�����Rz�f2��X�bh�l����L���6@��Ȇ�6�#��Jס<D.B��d[%���o'8݄�+Vb��-dv:cc!���Y�E"�R�mE^�D}]=Yh�1¶�vK,=if&E�GCc~��� I5����r3izz��{�ALLN���"'���.r�⽄����ZD�E���	�NX����=��!���o`��ʟ?`����g�^���"=���~\�m���q��I?y�d�z��y'�8rm'@�y]C~��s�h7F��:k�GV
z.�9 �+o�"�P�����2I����"��O��~��y�*���x6a��R�]©��E�((.��p3d��XQ��r�tL�dNZ(r�|(i�(�^��fb���ع�8�S��!�%�`r:��1���N���'�ػ�I���}����9�
cO�n��� =3��w�� >��?��nDL���_�Cp8��7m%V��P"��r�B��%+���#XI844D`�(;i�j,��E,������X�Q�'�;w���s��U�Z�U���<��џ���ٲefA V*�J�܊��ԓ�����l�^����������v���?m��JF���E ��I�k!,%Yi��4h����սh� �U�U9�sxJ�³�/ѻ��׀\������J���4E��D$�_�K��Ip#??
@�G���ߍGy���,����{M�+g�h(���Ε�_�o�,����|%h�����f��7�V��3�W����p���\�Ĺ�<FD/��\��D}�ڮ��#8��\�G�t�B-z�G�4�JK��d ) S �xI��1�{�ڎ���Jϡ���;�ǟxւ+u��Y��� ݖ��������#��_WW���\������9���������'�}#��L��J���L����c݆ud��hlj�5�l1�Cv�G���SϛQC���F�=��C������$��Jo_�-��ܹ{v�1���β�tET�~��3�chdO=�^Y���d��%��]��M�����,�}K[��L}������]�߉�Vn��������1<��9S���E��������S��l�i��1����	�����3Յ�8��.jK��7�`�'E˗���slt��Q
����n�������W�485�K�m��u������07�����&+�#(& Q�?(և���gZfE�>���Z�WڊQ��J�q��	��)����J�^b;G$R�<����j�����s�.^`�VS�V�=�x��Ф���h��U���<!!΢�Kz��%F"�)%�t|҇j��(����*���(����Cp	�)c�ҥX�z9C�hř3琗Wh:�Q������D��cT�I=^,NzΦ�&����:t�	������o��B�盷m����d����o>��8�@P:֔t�s�Y?$$���f!��(PLN̈́��'�q7OR����j��R�y��Z$D	 41��)�lL���4������1By�<T�ݔFxm�z

��s��{��q�hjl�@MQ۹2W����1���#UV�kU� �?8��u���b���2g��sˀ� �F��Y��d/.�O�S�� ����B�E�U+�3f��� M̠�w��B�Q#�"�R�}2V�O�&�B@=3���z�u�-XF��vԀ��#}����s���j�J5" u�%S��'Qaa֮]���n�2��6X�����ƍ�6o��=W�^�R�Bpr��\������֮!��bpp����2{L/���n��
2�E ��`K+����S�E�LII�ح�L���˳��*�Y�N�/+/�֭7b��Gڻ}x�)9L���]r|�&����k������z�g�ϾR��mU��m|.j��s&	�ri�9_@���@�z/�-ݣ�&�)�,S)/'���JK�-2�\b��Efe1츜����\��E�2�G2�T�u�_�rEG�;:�?u�/u H;1%W�Ǎ�!80�{�<|X��
EŹ��2d/%�+���4��>�sS\�O����.�c`؇�l�;�"e"Y�PxiCL�b���+�i����	2��_�������)A*�L|x	������z�LU @�`�8�blY��1�h�W�r�Kw�0��?�O�|�Dl��*(��#oy3J

PO���_�xQ]Y���2�(�����3d�^���?�ŋ�M��we�1ǀ�i-�űm�?T{�z}�D�"�f�hW^�[����i����@�X�Df��.֧P��{���R�����GוzE�t���ե���x�L�H�8�1�-��rt�9���͎('�ݛAQa.��ۅu�V������Lþ������WT�.{se�\�" ��D{żP�1��kQ��`�6�1Av"���LC{.Է`":�������8~��m 
��*�9�&�&�,hqWo?z��>'.@� Ejn3���=���G�����C��`��2E2���Ȁ\�� �)����]]r����,
�*�P��6���:�����j�������Cq9.1����?y�����v�D�������܄��fùq�zd��f�K˲���_RZ��",X0�����[�*r����娨*CzV*fx��I����ӄ㾪#2N-P�)� ��{K�젶�Hmo��U���Gk�\E����ZxRz��<Ŵ(�/�־Nl�����X`�P�k�@1��	g��"���e��]q�̕7B�r$山1S�]���b����v� ��E����/�EJr�K�$�56�S��r�OC��(O��a_� F}de�u���5v��{����,f�A�A(7��D�GY����˸���X�p�	���Dա�1<��~��|��#C�)k�J�D{g;zz{���wvuq�d]z	����0������MC��:p��e2�}��Ёؤ2�Lni����>���73 ���׭�����y�6().D���xK�+1� h���F0�6R|�o�@�pt�r���cf��{AN>]l����1N8^����u��'	~�+��߲���h�Sv����fS{Xx���}��e��#@�Z�j<��l^��1��i鿃d�ql�VTWW���ύ�u�b&ʓ͕��("#Z �(���R�]�b�=�����Y�?ـ���&H[	�c� �Z�x	
�3��يK玡��.���TV0���CHl%
�qIH�c`$��G����:��'#ޓL�Q����.L %2f��"-5�bn�x�G��'����}���D����¥|����|��p#Ν9�s����-��b�L���UQ��
� �R�!��BD �0<2����c4���śͶUAOL,�!�U�uI��V������0>6��y%xꉟ!�"�}?��T2�����>R"�]<��`�fݷD|�CQr���k�'� ;���� =]�� N��X�:��fWݔc�� ���P��7��]��"��	7ٯv���:� tJ馕c��qǻ(����Y��u��>ܲ�|��_F�'/����l��~���̕�Z�~C<Qĺe˗�^�r��j�U����~�z����������ꤛ�n��0Y�EP���Fbr�e����$��a[�oh�ĈWv��-����[yH02@��z	�1h�;�6�7�&�즧�	xA<��N�y�-�(//�[y7m݌�+W�z�Ӄ,XPm�����CII��r�_5�LV.��l����c�����މt���?�8E]�+7�|�?U��\�P��������K7F��j�*���#Z�E�#�h��LL!�:Q��0Agb�m���1�5��dh8@�r��wt��?��*F A�@O�Ǉ�������n�����
�{�W��e7�<��c���=��~�W��"�$��ǐ����OJ��)B��JW������&��;�����ZO �k�	�t���c���Jͮa�_��
��o��%�p�,<Y��dd8|�b��i�⻂+�pռbKx�@`���*��ؘ��=�{z�c^7!�����Xl��'���!/FE�%8+`pnN���w������(���{���pNN�`����G>���B�����C��η=��y�[�����OJ4���^.b��h|�����ʒ�J?�zzbƖ��yx<d{��cq�1&��&���q8����u���=�an�ifu��Yz�#�I���ջ�z�=���cG�]��](�U��W��W)����~��'��o?x��W��L��aY៤�-�5��9�@]E	b�C�i�Wg*ˊ�~%������3(�U:$e3
KOJ
�&�g������Y��Zx��5�-��i_$�*T���z��;e���@�~����)1Ud�u�H�ʚDzc��>?s8�d��V�w��
�eL�4Ÿ�J���3O��k��c�G��z챇-}�џ²X�ܒ��:o	{�(�6�e�#V?/���;c���H�q?��Q���"��3�>�cZ�$�̓�(��a\���ٖ�k���a�n����>�t���}�qD�He�ٺ��%���)�琽��C��h�_�b=����n=�7���_�@%��mfꎝ������J*�WP��Mg�+o��4@�M'	��������8�G'��<C_o?F��0�7�a������������MdV]�!���|��,�-�j{�$�"����c��D��������p�=w#��3e"d�@�	�b�1��)DƢ�;b	��	�T�>�Ϧ���Ï۵�2�b�C?;͘�%��J� `��>Z�8bq��N":9l���1�;���Db̮O��T�ҥ���x/�N�=�1���=Cf*�������\�]��T#gѨ�}�-��r�zww����q�R.A���;�DIi��&݉TT�;�1�@60u��qň��o���gPXMV�Gl�`@1=C�+�NS�n��&��$��3��%(�p���۸$��˲(²�U��L>ck��P����_RH��p�'���'���k�8�S��z���
5uN��ܩ����x�-{�3��\+��9�ӧ�X�Z��e1��񈁚���J��''C��v���\�	���	0I�ܝ6|�b��
�f @�6K񼻣�?�����U۶�����z~)�g //����!�M���@0hK@�ȫ�+и��<��Q���������zz;����zKf�C��,#SM���æ����F��;^�:^y�<��HGg��?վ����ʥ�u�wc�-;���Z:��}�2DZc�$�iɲ���N ����tQYJ{c	H����I:SU��'�(��[�ne=y#�t���O��'�b�����o��c�QP��8 �����fkS�,��YB�l}J��D�������pJW�&}\��V�<)�I�P����~LٳqLG�p��S��'�w�zMH�H��?8����Bm�
[�4���Oqݞ�v�o��4�~�9�����T5v폤����td6	���k����b�=�
*��"��P����O��'b&zK��J��M���(Y,���|,����͛li�3�<my��N�i��)�i��O0���:������ΝW�W��6�p�3�����{{p9X�nn��:���a�%�q�Zlذ��i#�J��X�?�D��$�֑�{�s��4����PuIFU��^[�h6����hni��l2��a�^u����ΑH#��hmmE~8%�%�f�`	H����y@:����fm����}qi�(��;�/���;R�����??���*�H�$0���I�A���)֑�xIO�ɠ����F����	��c����Y�刉�O.��LP��LlH_u��K��[�?���'�r�?v5��?��_U���V���wlظ٬5�|��[�;�65(����u(	v�[׵��ĉH�(�5�0GP�[$�����ߟ�\�7��щQ�tõ�CԵ(�U��fX�Σ��*��&��/C'%%��$Ξ=O�|�q��^��~+��O��&�N9����8��[�m�o��{���a�[.6��g���-m�v�:���=-�V��2�Νe�	.~��1Dz�d���CKT�+���СChj:g��a�b�&���=���~��mo��4u�N$Z �I�����l8Cۺh,J���.�%�svR�0E����~lڼ�����:kc��=�C�.��o�̬�uEx)pkV���H�2��Ī|�Adg�ʽ�Ԟ	�� ���&B�[��Z�6�3��Y�fku�B2Ay�&0�׎{�~5V6�2�-m��9߅/�HZK��+jq�-7�8߇���r��׿;v찭MԠ�|͚5�Jh��/o4Vl�������sx���d�0<�GP�$����<:�. N������	�O�b���ջ�w�j�����f�
��!�[� ����Bj('�z׻�������ڒf�lٌ�o��i�c�Q<��C��Ӹ�7�w݉��*��e&��Jlۗ#����9[�����駟��?��zO>��Q<��<���|O?�$�y�I���_�w�-me$6y5H�<Ɏ����h��$�f�W����Pՙ�1P9W�4\aG%f��+3SvI]rK���S'�h�UJҔVʒ�8�G?B��s�yR_��w��JL��0-P2RM�(~���Y�8�:���k\�̈�G�4.J4!�2fDV�4c� �)����tZ��|'��@o�~�� ��nK� �|z����C]M9��f
�>�Ӎ��Na�ƍ&�j{��@�"i����("��2ݳ��4���SOQ���}��C��U�w�]سk;j�+�v�J�t����=X�PO6�W4 2>B斉��z5Ú&�w�e���vHv�k�g��D^1_�b�ss(^�� E�G�btl���7�t��<S3{��̌����)��0�W�����T"i�X_���J�Yg��Ԫ�ZS﨩�6�]_W�e�h��|�-F�b�J,o\a�c~��EEY��|�g���F�X�+W���79ò�F�Uq�s`U����<�L�M0�J�&��R}�%��^N*y�����7N�E�#�$���ll�8|�<�z���o@*��ꎔ���H���Q�(�k�P�\J6�w(9'��ƥF)1_�́�DM���,�#��P���q��ٴ����T�)}�<��S�St�*/��W�@Q�c�C���`�Bjjkl�U{{�Y��-B��i�ɶ��Ȳ�B�F��b^Z����.�J���J��s�����W\�î�M�U*?��r�u,}���[ҙ5C#��W|��E�[fqkK���UV#''�,��$զ���o ��Y�����.Z�ڬl�MHEE���*�ޞ^���ݳ��^������\�mW]�];wa�#��f7�x7Y�.����o��JJ :�%�@���Y�*mWEeş��%���@�[i5���ڊp8��Q�:��,��q�[r?gG�f)I��Dht.&R�Zp�Q@J��:s�)i�/d�TD��x3�Rt��C�*͌i������B	h���ʌh<.�`c�Q�-"�$O���qw���"#�P/�i��H<�]���i����i�T���8@ڏ^�5�(��bq6�D&0�����*g�wҞL��d�ף�0ߘ��f�x���Y��ǢĵHeO����ˇ�&_8��X|yd�b���3{--mX�l9��!<p��۴q�����EWW�x�)2�~�P2��$�ě�&l�ֶ�kK&���֨�F&�T7n,R[#������e��ã8�t_��W���?��G���|3>�N�c~Zp��1<���>K�L�p�6ӓ�VM�i"�駟��>�1�9{�\s�1i�-�ج:'Q}�%��^��DM0ke��&��j.`�N~�:�A1[K�1E����}�:���Fd���HD�2���TzY���0�aͤ��1K>d���9K���L�hN=�B³�Ks��55�g���c��o�m�L2'v��P����C��"�v�^��މ�?&��'���1{�ݼyy��f�5vi	b^ZȦ�5PTT������s��Ç�䏰rU������ĺ5��w��j�	��jfm����~�@x �����yL��B�~����W��p� +�Ybu�������:���~Ѭ%�������׿n�����G>�a��G��?�!�?�_P�'� N��Ҷ8ɵm���hMu�M��8LrJ��53��o���l��ӊP�a�3���1Ju4ڷ_ҁ:1�X4jl���}K���۔ʘV8i�jN�G�߂��w�-�$���٢uY>�D�ܒ�y;�z��6���S��F��L��yO��n��W0�F��4H+)&'ra{����i/�׌���.{]��:і�@�ѻ������L(���6�Ӥ��b5l�I�U�]{�஻�2sv�����7��9ƣ�&1G1R�����7�Ϳ���mo���V]da12`�Ôb q@��yH��6&�I���N�8���,��f�����˗�x�v�<��!9rʖ�ʲ���y��0��PF�9��_���:�'p�LG�������x��q��9hG���A\h��q��9�9߆֎>����F12��h$iZ	��˰a�N\���Wc�57aێ��m�5ر�Z��}-݈֬����+�y��p�-���W��핯ƪ�kmmKk��yIQgeV�$�/�%��qb���ld����S29e�{��.3{fRN3�����R�1|c�Z�ɧ����x�}������q�y/r�'��R�q=1��D�γ(VKoQ���3�JI�+�4��%�	<5�'������R�19>1��Q�@;����)�<��3����(�7�kuu��u�!�{�����N�:e���Si�S�0�p�	~��qr
QVQ�R�e�ף���P	���_�k6�~�Z�c�ա���u�ylDy����kQ\Z�"�P^	�fd;6@��Gr:1JعLv~�@ol��Hr����b���Q��X��qɢVkk���*�2�'���/�%�rp�(�jF,p�e���M��G:k����j�4������T�U�$`5����W��lM�S�������-���<���$�lfj�7��y�0EY�@:�d<�9"���5�?O�`Ö��b=u+��]�R`&�{zN�����_ė��U|�{�D�,�W�֢~Y��pi{M��은X�	��@&+�+���-f*�wn��d�%�v(Ug��LM��=��Ȟ�	�L��@6���=��;e��eD�#����3(�O�Xh�LJ3� ��x
㑘��b���I2�)���O[:Э��x<w��jYm,�	���1��w��E2ܶ.����Ƕ���UE�(*)%�χvku�.�Knɽ\� �`�mW�* �܅�h����)+?ɐQ_�+u��V�+�F��xO�0az®�KzeH�4�:��@5�t�ys
�7�]���`Ҹ��p=��Ӑ�3���/}���җ��<�0|�!:t���$y,�R�l6|����U�U�kV��o���?�����7��X�,��p����S&����
�e�f�ń�D�m[�b��U�ή�N�$7�(A[Z�CV�^i��w&"�IK�>�\*��>�Y�s&�3�\u2��w��)��8�o�Vi�� |̋ۙ AP��!}���@{.I�".��� d9\CYz״.d>p�P9�d����v��`%��d�3L���B~U!�'c�R)�$�%��^VN���6�a�q�I�?C�S;��i�<#(�Q("SM��gU�@H.�k��y�*�&k�f�=F�	��۹K���v��흦�9���
�'��;�9�H����<���~M�{��G�ܾ�dR��n����&���^8/ϼ��;ׄQ2���B�]�� �G��Q������x���o�>��W]Y������ℭ����ج~_���ɺ��e	�X�~��sj�ז��$�˧��f;qR��.�ڌN{�k:my-U4���im~N����eOND������H1m=k:��.��'׶���_�Ό�'4ġq�Yh�=��|�K�ݯ1ti�5�e{?1P��ˎ��V8^�YrK���T%֫�y�� S�P#�#v�����<}`�6F��]�6���#�6o�ޮ�9T5P�`u��`j������3f�ة�|
4�D T��1IMr��),,"�����\���V��g�~Ɩ��2���<==G&'�I��}MD���ⳟ���w��o{���w���{/��𶷾�|�+���݇?��?�o���o�V{)?>~�	����A�ˆl�����$���U��9S^*S�fʽ��A{<i���X�X%-A�9<4Bf;ayV����h~'����ʪt(�Ը��ĤM���tj�|U����g�%���0b��DO�69%c�J���w�*m��x1Y���N��w�P�U�%��^&N )<S��0��ڛ�V������
�r��>I�ـ@�Q�����a4��R��C��y1Q	��)�[⽀ҁ�E��α��������:�)��V[�.4G�buz��yz;]��;�Zv�9Ŧ��W�ZK��cT2�bZW��,d�3��U��(-���lt����Ǟ����PMQ~ժ�8�JK���?�	�����h�����튵%��x>���5d{AD�);j��ɰ|h���Z�/f�|i��sJW��:�x��N����XB�v��n��D�ֶKK@�����ٙos3�d�ez}�VH�w�S��}���CП͎���Ƹ��2��7��}S|^k�3��UA~��jg������Z�,�{9a��*U-m�۔�T�a2:�~j����j
���}��3h�DvN12���j43�d�c�"�ki� ����$ź2�̌�]
S	��X��RPu��@p�ؕ���A� DA����Y��n����s'�ח?� �韠���j�4�ڬ�oX���P����$�,+W��g c�n�)m�|�(YiG'��fJ�}�c��Z'>���r\�}�lۉ��:l�q�|ͫ�y�>7�p�x͝w���x'������b�Gc�qh���j�N&��ы�-�����6�� �2��|~�s��S����KZ7m4��a<���AhV_3���,]V�"P�q�(���)���Yv�e+�23�A�|���䈔d���%G'�y=f���2������l�`�o:������y~��Udb�l;���<�z������Yc��h�j����gC�$��Ity�ڜ3 �P�����.\��j��kA�@��"i.Q;ɸ�c��מ=�Ȩ��Iő�>Vd��$c���T\Ƌ՘S�B����^�n����W���[,�����=q�k_�F��]��W�����cO#� �фxl�_w5�k��HI_�|�a�˿�;�z��������&<��ط��oj��~�?~
�m����:�l����T���jӖ���f�g(��`���Q^^�3g/�3��Zڻ0�x�*�P^]�H4�N�ѥe�O�	4�����!|��2�?�����U+144���J��:�+�O���#d�!���sK$�*~`�țX Pk(��(��N娭@�>��?�o�#@y��9F!��'؁�v-�]�8�шm(��ތ����n�L|l���g��Ӊ���hi>�ޞvۻ�W�n��r���A����-�%���y����ʉ�-�Ґa��<�\�յ�.���$vr6��H�HC-��s3R+�Ck�1c#Gbr� 9A1���l2H�17�e���do����Z�-�j�%��l�,U�Y=��� ��Բ�����3Z"�u��};�Ց�2��I���5��}�6Г^�A��;l�� Y������j���[Z�?0����8{�,:ot�V�ۘ��8�"}3N�:���~L�e��lu|r��tv�څ�嫰e��-[i3�Y���SO�3]Ӷ��בc�p��I\�Hp�3�%��dz{�q��~<��8{�4��5�Ud���X�fn��&[:��ڍg�z��d��#_��k����3'�L�I��X��F2U-2(.�J���K���Y���s6<!s}}��ÊX����WC	
3`{q���r�XQQ�t� i��ڳg7v�ډݻw������-���`�D�ǫxKn��?w�r�4x:g����{:�Z�(��a����l�H�;1�����������UT#�_��� ��!dP�&#%�!��ɢzr�������(&�Q���gӰ����Ij6����N��I�%�7aS�!9>���=����?��=�S�~-�o����3ՙHL�~��ػ}�$�����>�o}�;dP-��.�8���2Gm+��b�IG�L�LQc�y�����E�K0Iv��9�����x��os�Do���'O6����?���Sf�82>j�rdl�yJ�����[] �8�5�3��)+-!S��4̑"���~�7���*�=���{���<��CK�77/lFT4�c���S2�NA[9kbHc�yy�C�`&���U�6�M�r� �}�{�p��GFH4�e��|�8�,Pi[[*�/�r�
f7��PD@��3���?n�`ҟu�wQ�]rK���4� 5<�@qa�IR����-[M�懝�Ώv3Rm�6���G��7p�� ʖ-��1:ډ�XB��Eޭh�F5�Y�3�O N ��H����@��G{w/F#1���"�C�
�x���&c��8���G3Y����ǡgt@�{ah�@�-��w����ƕ�Y&�h�p
�����m7� ���x#�����T�dRN���1�' �خ]A��d�9y�\t�w�S_��x��!�}�|��x��ވ���p��p�H;��?�Ħ����ˌ�(���7B�0���4c.�"���+�ϟq�l���FQ\T�;�x������������� �ε��	Z>?;���:�C�Hi�z�aks/�pJ]�����6�2d��|i7H[A���z�Y����b�p�ղ���*�����DV�XeZcL_uU��508��[�`�,_�Kׯ_k㻂̋|�̙3�JLZK@��^6n��Fj�A$�1G�S�/55��nK�/u?!�&x�I�o�����A�����09܆��VR��LQ����"�4F�z��݊��!�V��fËc��KJ�E�����f���-m����(� '��4���K��̗�g�3 }�@�o���wm�H�<Є�����5�L��}O��o�oӝ(�s�DԵ�IeG�ɂr^Z&u�ːd��^���g{���+��k���X?�6C���X���i�#/F_W/�K�и���B��-�я��!#'Љ�ي%�C�R�fbº �*C'C%�YlN��>�����>�%l��j��#;2���VvCH�'m�i2�2����,����Yv���Yv��BI�6;�o�[���^�j�0/�3g�پV1���n���c�?����|�C|�-��mWY|:y�mt�-��?x��I%����47�ܹsƺ���-�[rK���{�.�6���R���3H���s��l߱�ډ�����ԠE��j�(��Z�lb�"s֮����뱼�ӓ�;qG�C��s�L�Q[V�-���W��}w݆=���YL�F�͠��[[YB�Hp�I�z����8��G�c-^��
t�8�]V�6YlҊ��P�"y:;��|�c�[>6�0�z����R/���<���]�J��V@%��@�u��Vl�?�Zz���/�G����O �W��׾�����#6T!�+�[X �}(��0?�y�P\�ca�1�>���#����f��h�lʖ����,j�ʱf�r��$�6������X���b~)V�\�իPZ\`����Yw�0��j�S�e1�Ņf����>f:���<zY����z�sٻL<��������M$ḅV`͚����h���rҗ��ɴջ/��{�8��T��l����k�$D�����?a����O⌑�z����_GsW%ک�̳,?��\�ڢ����c�Eey{=*��̤Ȫ�Oۙ/�lb�w��b[�Y���a�tt� 9��Ԝ�|>��� Em)qgg�"/���x/^x��H���1R2U��ǎ�O����Ǎ7��?���.4T��� �)Y �e�"�F)�1�Y$b�� J���J�)��X;�����5<��o@-�f,1��#��(`�盢�O�L�(Eݎ���M6!���G��+%.M�~����Z�%�ؚY1�=��X�n�3j��_�������w�aE#�ݷ'NG<C��z�ݻ��ׅ���fQJ����>��j�ه0��盵�#?11i۝���o�������V��~ޫ������TϚ^��u/Pd�^Mb�����J��g\rs8y�M��i%�U�ŵu�-���3�w�{[��i}�������(.)�UW]e�U<��-��ܞM���(9Kv��-5�JpՆX�����<t�����G[�l����<;5K�La��34"TO2QŨ���1�Ύ.�HY�x�b�4R���\���w�ID�a������h��$��Zmtt����y��{�5���	�'F�v�����tK�&~jLR�^k�m\r��g�mrJ�@��G-�T��sd
l�ylL��G�/d@�y
 d�$'�&0�� c���<{�$�=�f��݁3�O�v#Z&*�~������5�v�<A :��D|� {�1�ʛ߂��2����]���*lڴɬ�Kq_z��E�g�4Q<O"�����K�_N����ഔ����=6U_߀��<��8}����r𡽭˶�6	U:z-�8��VK���*���kyY��5����������[rK�e㈆^�n�T�x�k��"�t�ж���C?��Y�C��1���h�G}CV�ZF �G�G�@Ws+źe�z6Zr�T�H��3P����yj�`�m복N��a�?xm�d�E���w0���,��El�Y����(g!6֍sǟ�>�q\�g��f�s)����[��~�7��=��N��l���z�jJ����b��SK#��=76�ވ^ʹ�n��@�ֳge�I��o>���[QPJ��K������]:��H%�� ����L2��i�EGG�����R�����r�%�i9�:L6�u��1R���t��hlO=�n��U�Bp{�����>���׬[C �Ŋ����ڌ/}��6��G����6 ��-�`�Ԕ�Q!;�˳J#�T�ܾ}�n݆ё1|�[�±��lGE�*�F3�d���nG�x,ƴ;/�mn'����"S}Җ�7�p�p����U(U�%,]r/���������*�~;�_DK[�~���8����r�H��8~���}��.�1���<���G_G'6�Y��{� |�N#�`Q��
d#��${�RAg(`��� �\�M�Ţ\��bP�i֚n���f�<C�j<���.���נ�����f�enx<��?����c�G�z�W߂�ށ��B�{������@[`��<H�a�l�g~^x~��V,)����'�Q�=�<����f �M-a� C�&�&LQ=�@�Ӓ��9�0��*�_�()�'[�v�e(/� ���q��**ʷ�#�	F����F��,��`	���Z�;mx���y�%Kdw5����ŋ��{!C&�|fX:2�o��ɘ�:A�v���~�mK�5��bs;x����D�,�O�(^GI&g��!�0)I#2�1RU�,�����5�\�t̾����\W������p-����2��e��"��b[��=�á\�#��S�p�ׯ�LS7�l�؃�b?�y���g�pۍ�"������`���O���� �o&�l����e��]:��e��b<�����׾Gѻ��ƓSRԔJ�,3��5��\�^\8} _�¿��]���ⲯ�6�#gz����d��L7���	����y#A�HL��f45]0���+�9��N��ٺYG�h�^��s���V�f&ۙ�$;���
{�3�2��"L���S�d����L��7N�^�޾~�Њ#�̳�d�L����)�*V*�μ|-�`>�x��sԶMf�~�l���-;91���m[u2����h|Z��Ҹ�8�*��d=]6tM�J9���os(=�<b���ւ�T�,U�b���0Sx���l����b>a�?��l%�r_rK���~4#u�-)N�Ej���B;h,~�G9���D�������V�ر���F�l���+����߉��n;u��Ρ��6��Y6ZM
�ѩJ\U�ITQQ9֭ߌ��:����&1�A/A�O��I H`||������S�	����n56(c"�O��g��]��mlںӔ�ۛO�/?�{��U�cx��}x䱧p���d��ƌ���0#� $Y8�D�6����6�D0���������F�9�,ǌȘ�,;�d,N6��A�(�q�ڱ���
�����a�L�Sc���-$�O%��=���enO�U+++���a"wVv��_����~���nY����LD)������M�ixRJ�lU�Z���% �3~�眳��1 ������{4�������q0�qY���^U^�!�R}>2Z~S;	��i40�_�[~�����IO=�8�˰!�ں�%��~�����[D�U� U�۶nECC����Q.S)U����Y�z�D���9��Oģ��(5v��=?}P"=bvV�`C?+H�6�#����f�dMI�wiE)y�k�#fv�q�R�xO��f��QlϖYЃdN�WI�?|�}g�g�SL��`/bd��%%غi��܁뮹����b�RW]���j�ޱ��x#���j���[���|e	r�S��Z^D��$K�!�EI�yĦ\���"7����8Yp������l�IKP5ѵr�J�Y��y��$ �&xvtv���|����w��O}��8t�(����dEU�#����{���޵`r�*�L�X��V>�xb�y��y/�^���,�ev.�)��P���	�Lw^1|V�'��@�^�C�����,�Í��0�}����J�H,�?��Ua2�����u\6p���/�S�5"B'r!CM���$]"�?��1R�F)�>踙���.ú����d~g06<b�2l"`��P��!�@��?�3}Y�4��R���#�x������U�.� ����_A^.�����n�]w�˗�8%�g[�������z�z�;Ex �_��V� �@UU-6�ۄիV�z��-[qs�-X޸[7o��߆�n�	�6l�����s�Nh/���Dc3���(���Mٞ�	E�)����3S	�Pď���
w��U��)�=`|d��׬�u�]o{��ڞLY())�}��W_s��24-C	�����O>���^<���d�yl�C�+=U��@.�Jl��.vL�V�H��6)�l�9?�ͼ�\j`$�fLDC��~�m�m�@Re��+�A第�+�����ᷔփ��&������;^mƭ�nVKJ��IBܒh��^�k��,��f�R�z�u-��-�/��Q��K�bkB"��;�gAKJ
	0�6.J�C^�֫�566"���f���}�~��)z"��,ZU�Ƨ5�m�b��PYi>Y)�%�T�8����۰�c�I��b����s��Ȅ�NQiÑ��rN-��˱~�Zc�9L��L3mY�%#^�z5�I��FFl����0���Ҍ֋M�gO�Po;�HAC>��"2܇҂��W���`��	�1[m���O���}֣i�S��h���OK��R�e����-�ކ�B1�Z�;ׁ��ػ�����s:�Aqc�"��`�%���L6I��K\�.��E�ʲ�&�TY`�!fm?"u(�6��D_&6�iP
De����ߙ��S<.~�����~_�6&�mC"b��B�עU�%]r�8΁����-�>�id"�����3?�3 �f�K�RlOADs�F���/�� ;g�Wd�Nf�4�.q���,���;ś� aB�Y��l��C#c����H9K�H�f1=�VO`���!� �̄>���C��C� ,`�"��vvc͊ը.�D Ç����&ua2�ҲēQ�>{M�ϱ�fx��y�&��ű�����x�:�Z(�����݉�������;o�������z?^{��زi��+�����o�7~�װ}�F����������ƩS'(�Sd�#=����( s��,e��`2B�J���#�v��<�)>L%�d�.�1E0�h��ՄV �`rs���N��ד
V�}X�O�,L�	t˕�|M�1�iDh�S�M(3�d���f�����k�&m�Nh�2O��gfh	k��eÀ�����d1Bms��f��o��N���|d�|F�w�-���s5Q#���/��_n�$y>-�r�"pb|�|B4N�����zn�Z�3c# `!������k�hf���e"uX,2��賵�Sd%�%3��0Gdr1����O�mCGɂd-�L\���168���	$��`����qD��̀I�?@������x��&������:��!_�a����f�5A������YW_��֡���V9�E�E6�;C������4��z������z;����p�5;q�M���W߆��r�a��Ξ��݌GY�(&c�o�痙Cyi	���`������@ey1�0���τ�&q�d�2B"��N�1Ĳ�`�α�M_Uz��2�s�IFcG��e��&xe�F)EzI2�77���CS�z���*�|3<��������Ty�*���#�H/��{`����=(��,;�X"FP�P���4�]�^]rK�������ȃȄy����ڂv�H�c��l�SML����S��x�g�"�42�����m��y�(*)�����S�<*����d��j�ZED�b I����1����ǑC�PTPjlt�ah��VI�\���Yx�Qj,O�T�4v!���\N���C���h.
�p�i)����M-�s��ڲe����p��)��*�RH�V�\���B3�12:J �����1����^R��lb��?�)<���f�T�h(���6ld8�('�o޼5�58u��)�+NY�������zjI䁦��ΙǠV[)��Y洙�)~��ál2s��ay��x�`�g�`-��Yvv��|7��{�Z�����B�f����ܬ��OA���>�:SL����䷙���P/Ξ=��7�'�xgΐ��C��̾K{��,�%��w��O �n{�Z6*�h�@�q����1�)1��"�&�<[��q��^c��֬E(�g�����#l̙ó�6K�4M�gB�(,(f�atx��^DOW?���ϐ�5�߅�ɖ���L��n�ׁ'eJ�1p���iG�ؤ�_�&5�k�co�#�*))1�0��yz3����rS���O��V�h'Q����p�]`����c�����IJO��i6^�
LeAFiҚ�6�̟�-�y�EŶ�^�5773�s�z��\��;KQ<�S1c�y�>����3��p&���"�s��ك��#�Dl�T��L'&��MR\w~���1��L�ҕ%�
te�;� ����ǆY��l�>ËFG�:����h���ϳ������4:l�i�-�_Ǧg��J,NZS$uZ}�M4=c&/�]��ͦ�f�AV���al2���^E�((�BQy�cI�^�����p��I6X�F%����hd"N&׊������Ϙ�LII��GJA��Ф�T4A�a����x�*�Y�x_��X��o ����Pt�؝{U�A��]{�tI�u��>�^g,N� �Y�Y�X�,��!+����׾o|�q�7(7����Eo�`΀򤭩���իWcǎ]f(����Lz
��˰\�[a�@0D1�����n}�F�SQ�4�BY�1��4�"3LME�$��V�2�v�Θ�1�Y��,�OC `s�'1;5���@u��0�C(gcÚ�ٹ	۷�ņ��ظn9�m^��ee((�Fq��66�v�����ĭ7_�w��M��?�]�և�O�3��I�	ż�1�7-�%��4�$B����4ɴkZ�7H��G9S�ʦ�a�p�4R���$Y����;���v��z��QÃ���0ۗ���,Zۺp������a �I���)���)�s	h����U�j�C�ݥ�4�=�}�j�����{����M�u���wn�ؾ}3'���Y(+�$t�&������9���j8!f�y��1��w`��]hl\n����e�EŅd_+�Rґ#Gh�f;;;����c�Ao��vc��<�,^q�ͨ����dYi3Y��}�~�93:�|�
c�'O�2	R��F{���"S��BE��L�L+�����)����m��k�V�YوUd�֮��a�j�^ӈ͛�7c��5ؼi=6m @��z>�n�
�Y��V4`��Z��[�����{��ـe˪�q�*汐�:����]�*3���ر}+n��f�T��	vDn�W����n?~���ܒ�EpF�<���T��ȯ!GIВn��g��#rrV��Gヲ��o��lf �#�8|�N5waƟ���[�|�VW7 T\�@A)f�s0��E���,R2��C^I�1�(��u�aj���?(>�ʠ��TyE<����"t�1<)�le�H��T��A�d�����3P3ўN��=�FF$jÔiGGG1<<BzN�� pڹWĞ�}S��elY����/#����|f#Ã�Q��� �Ҍ����"/��Q�@_�JKm�U "���X�(g��m�g�a�^nl|܌������ ��;��z�Z(B��6�=�y;�W�kw�޻�����[񎷽	���N���o~�=x˛^�����x�;ߊ���;�����ǣ�����.|��7��n|���}gEC?t� ��u+�H��H���W�ى=����`I�kj^ډT�QO%�xᢍ�˪���α#������ܒ{�;a�Ԟ��}�RO��S��]%^j����h�H�����!+��x*}�x��9<�����,'S�ՠj�ԭ\�뷠�~�YH�e!\R���d�`,:e[kS9dl����l,���|�6_+�CaQ��[*�F����=6�h{����Rn{[��wN�"���h?@���H@lTvHc�8��+�l>P�񼮶7��&3(fX_W�_{ǯ�[o�8�$���Fj�]z�������'��֎@[>�<y�,��x�+̴�D���Rj�X�gU^C�H�k^�G�#}XG���w���7ߏ����(:�/�� D�����sg�����@o.�;�<��<��/���#q���?w�΢��<Z/�#�=c��)����q����S@N0�?�;��1Zve8y�0�?�M�N��:���,��zmX'��avT�E@c��*���/���$�ڡ�ݰ����(pU[�%����r�wx�3�~��z&���s�� �_��S�@�� �`���>5!c����1B1y(C� zߐ�֮~���DI֒����2�,;�m�Kz���P��qQ���5�D}��He��z������4��*���k����d���3hk�¶�vR,-AWW�05`,���fk������ڪ���f�]�p�8~Cd��kc<�����TWU��C���"�4Ya�]��֮�2�F�c	���S�>H��˰{�.Y�v"���m6'��	���ً�۷�e�M��أ� ����k�0�J�d�b����g~8�&�4��,\�
�D�l�9zĆ*N�>m�(�gxzN��P�l����3R���ܵ۬P�����o��n��5�x/�4,��QQ^I�~9J�KMӠ�����S@*#1Z9��
�����[��V]G��5�1�#`ն<!�C"="���ݼa��I:qs>��9��Q$�ʢ�&�!#�Z��;0B��E3��"�y6���h����.�nGA5AQu.K,�gLTb���. ��59AF���8Y���b�v�����־�G��a�N�iǱgP]��tFW.�7c!�
���9�0�nێ��"<��sط_:�Y�Qԓhkb2�����ta8r�Z�[��ۋ�d�G�6��ǎ0�y�a�;w��	�=�"�
��@5f�dڢXF��5VLƭ�G�-O�N��}�d�����f�y<2�]�v`�NY���q�O<a�7�z+V11t;h����˖��؉>tn8��+V`�pyy��klBKc��&��ذ˖����b�_��&�����z���d�~�y[���"������X��5�� ��}�����!�
ګI:�iA��ܒ�q��=	�@U�ջNIQ`'�o�O���!ǅ1�,��G$Hw�G�&�2��� S)ݔ6j�?Fb3ZZ�M����&�H��5�=��	21�Tb4	: 峲��mH4&��Yt��Z�Hp�����y��O�jL����ʸɒ��#'.b����%��%i#iiQ������%n{�˴�?e,d��7gm�I*QڪY�^dYI3�zN*ZB[S�2��-�5��O`Pj�{Aa	���FlڼŖy*M�2h}��92���E�ؤ�y�&����o�!|��dٍ��N[ݻw¹!��?���)�2VUu-r�
l{�,�p���WC TVաq9��lY�KW�^�u6a���ظq֮ۈ���`ٲF�%�H_Q)s��X��o=��'O�\S3�����iKK��:0����ۏG}�*�2.��3��^�ʋ�|�j��.�_'8�,�i>E���ebOC��	�̌������ǿ�$|��Tc29���ź)�B�{*���|��JD��*�B�F���tO����%$�������Ȯ���E��F�Mf&tņ�r�<��}�c�*��E�Y���s_{���;v]c�g�F�G��l�Ԉ�����%��+�m�6S���fQa�M�8q�T��������r*�6�����#�$Hj�,3Kp�c�f1�*#��N�Jt?}�,z�cz����Ya�؛�������뮵=�5�PN nl\���,���딽���f�������1ܧ��'���-F�^�[�l�ب�G;��nĖM1�<i�R"^A�uv�1���5)ĞAFc�E��'�ى�˲M<���G0HV��b�Q2g-2C��Y������1�R��$��=�{�~-������:!�=	6�[;��/�.�_7G�R�i�546��c(G��,���sG:	��c*P�`1�tJ@J�F�&�ͥ�_�p�M����Nǐ�8�Gni�D�lbK�0�M���,���L���+�T�/��}��o��-M���O}���e�F���g�ѿ�8V���_L�x��z�j��8�퓟Ǘ��3T,�VlTc����$��SqJ�S�Gư�F���Q]FF���J��_�U��[�1V��&Yc3�������_��*[�$�Z����J���QZZbƔ�@X+���&�=Ɔ�+�q��i|�������+������g�?���L�udt��1l?�jjQE�}:�4`�̹3�H� �!��&�j�Ii��gգ
�ԫR�/QH�h��f�5��и2
��Y�Ȯ��^��{�i}>@ f{{{���έꀖ�
p���ܒ�Ewj#")j�f��"�;v�$I+�� ��j��kϟ8�Y�D�0��3Z�23�v�W�&d�d���ɿ����A��Zh���d7Re�
��F]��J���0��<�H���>�wϝ�*+��/5(A�G/��B8���W�۷�t-j*��;�M�=�t�&Z�R�ղQ5!#KL�.�ym ����
���V3������>���å�D�,��L�Rک�l:rG���l����sZp��i�4_�e��3U����&p�𼹥�6Ը����L_�Y�޺m>M����{��
PFY~�#���,��ڻ�'��ه��A4kL�B+.�t��_liGo�0�F0<!8jӿLF~A	Yn=֭�B[B�����=�x��I#��5-��
-m(h;���S	�co}˯���gy�����\R��fݹ*Ē[r�Nc�8?��H4bC�!1R!�s���l�/�8�9in�̮͐�
H)�촨_��ܑ�����5���L�"X���^M�ɀSw��(�S3Hss|��M� �Ҋ�B�{H�='O5��������[o�޶b�ʾ�R�7��N�����&�n�zlܸ�,����;v����z<�L� �CbjE�c瞽͋lk���]�#8~�,����͢�b��5ƨ����|�ظ�7��ʶ&��j�r�*[b�����W��ڽ@t����a��^�#+�OX"��L��a2�=�T��DU8\@\���Zv*�6t��V�ԣ��%�((,En��L������i�DN(�b=;�шt��e�����O��W�?b�b�CC�ƌcd�##��6A6=����L�i���v�#����/�s�؆"�J%yI��ts/�}���F�����w�<>TZ��la�&(N"�hV=5M��"������0�����&$<:u���f�d�/���x�?YsS(ga���.�?��y�2����|��>�>���a-��Ρ�f����^���)^�cl<������DBl��H(Cq�j[9�YNLN�jп}�~<��)�����(7�r�� �D[��Ƣ8u�4��zym�%���N�:��|�W�c C@��*�����|M^IA?�g�J���U֒&(��:Uݲ*�h�����>�e��8A��2��E�%�ڻI*P��%L���Ǫ�9A�{c�)�^��z�_�����i��,V��Em�-����L5��%լ�S�	�#�e���(��A�ٽ��E8��~���c�����<�Rc��X��
�I+Kn���;��Ȟ���Taa�l�mny�h��4#�HFz�$F� �P�[��&*d�Le�lMco�"�R���6	�p� +De����?�g��U��y�@�=�	�0����_�ZT��+D�l"�ɦ<��T�5"�,L+V�^������qLY!���u��)>z&>��i�,�"�2	v=�/ 
�]f��6�F�Qݸ��4�Z;�������s�O�g`�����������������P^�g�u�jPQQ
m]\D�Z�m�B����Q�g�k+PK�Z�g��ٖ��:���!��4s��C�9G�;ś�O�&�5luXQY���N��FI~��V]��eG��asN!(��dq�dr�T�2nG�dDz.�Oq?h��7�՛��^��U���·pם��Rj\�"R��5+�K��&��I�����͖ܒ��w�ƶ�m��z赕PUu��.��n�����zq����JTdC	fD���k�(�b��ıD�Ly�"&Hf��I�)���X�E�g</�D)�V���14�E0�;��F����U�޺ɦ������q�fIz��0IЖh	 	2Ϙ�H�jK
ދD4�����Q��I����'�s�L�O�R\�s^����+�F���b��| ����KPT���mA���B�\������b�ޫ(F�a1C�M;�����H6�y�*/W��O#�S1I �O��?��-��d�~D�������PK��y�G�@��of���T�:U�!�k�3�B��#�b���d�3�IC1�y�_�d��8lNn;�Op.�*g�9�������6o\nU���� Ӗ
h���`�%e0��)A�C^rK��͑��-�N;�EW,_���݅z�1C�^��?x���K�C����JD�d7�D'�����{N3���U0�8z��s3�y��HҺ�s�]2Jo\�.�
HgP��C[�v����<VT�92��{��'����뗰a���Y���^t��R��C]u�
s�6�}���"��)�� 4�'C)��K)�O#cc�JS�0��WA[k���G3��?��iP��{ZSNP��AU�̢��	w��Fܸw��>dh�V2�4�l&Y�!TR�W�=}=����V���E���W��J�W�a�J���
KYЌy��)��)�yOAFN4 .����������[����"`�~��9���5P�Xij���o�o�Moh�ja�t2���<�w����Cx��ob��Fv��/ۏvM������
�6��MI5D����Z�+,�%���_N�V��$!\���8��)�@z���"P�9EU'�K2dQ��4�ɬ&�\�j�2����5n�<��z�Zi�ٖ�|Y �Ǥr�i����l����9,�${��bx~��������翍�[�F~q���LR�� 2B?:���0�!V��i��0٤�b`��%(&�͐�%�S6�
�;����3�T�����)k;d������ Fzۑ����u�mo��@�u@{��ƚu�|�J�(}�qw�i4�������&�>��(��5�̱��� X��R_���&xw�b�/��)�k�D���x��߀�)��Ҟ��x����+,a^s؁�'�\���a�%i��I@��E!�u^@g�i<��w���̤�ζ6t��1י�C�1#u$3Ӳ��I�% ]r�\�)�CR�M�pÍ����e���gN����C7B �N�@�4"��J��)����n"��-d�h
DP�O=-g�P��3̈́H3gP������1�}|�h�$��		�����M|�S_Æ�7!��
#C#�ec�<��Y�E(���
@�*m,�&2LQԆ(�l���ض��#|\��3�h� X���ڪD��"d�Zݠ=��q2�@�;Z0��� Ǟ�3I\�g>���c�u(���/�g�ۇ�}��x��������L���7�v3&�Q3�'�\F1Z������ �����ڵ����p��	�?w�+��.�b�#�C�!��-_���������8�Jl�A�_*� ��M�
�46Bf� ��3��M�i�S�~�U��5��06&C�5u(�:Zm��-��.�%���$��6,�Q�Az�7�xr��r@�ȳ���x?��*!��g�D��)�9c�b�R�$���\�`�TN��N��R��" e#,g���	��H?���0�$�e'���ݏO|�hذ9妏){��4|~��#h^�b��q����bxR
�j�itr���g�	�Y����s�}�A�سf�5��w	�گJlNy��zR������Fd���x5n��Zl����%�`�d~��y|�_����Q\T�={�ō�8;v/�?<��Y|��_DOo�c�qOc��mx˛��c�������7PW_�w���PT����q��3��(��AYu����?~�8v�4Jx-�,WC3^��K ��V����E�>t��Ed��>� �JsmW��MM��5�U-R����m5��:b@���%��~��A�	K$�
HE�d�-��û@�΄7 D��C@�%�_z,���O�r�.C�N������;�{���e��攖��2�!Q[��5��x:����M���OF12�wǱ	[Kn��٦���>,�&��]��2�6��j��Q�
)>�?��`��|_���X��啳�$��?�|��b�{�ַ�W�l4�J&f��S��jٽ{W����G �&Xv���������Cں~%J�
ϟ<���V�ݱ����cώ�dE�*�ٵw�~�*K�JL��U%6��fE-*J��226b� ��*,M�%�ӈK�,srb�Vc�8�mGKoC!�(4� U,}�qI�L�#ZP��r6|�Ί�;����/�cն�`��~��WڹK|F�E{\pR�K�AhLT�L�����cj�5{v�{FT���c�j�~����mk���̑�`2٠3|d�_[kK`�؎�Tq^�堈�����[&�G��}<J���`�1NM�(^�@:J����
�bn^�1�,�z�eJ��6U���PRQ�{�p7�+�.��Q	�DLK}I9ݾsv�݉Db�Ν��(�-��++"�m�E���a�r�}�mX�P	�oL�Mab4n��XW�d4�&��)v �Ȉ�,�J��St��p腃�8���)~3��Y�yT��V\c�!se9Zy)����M�EZ�!+8�d�@6�0��-�%����uz1�ʿ�Ig���+]x�ZZzT@)1_3��V;�|�"�]��ib�
��k����}1���jH�"�<�eQ�l�`�]v��M��1k���_��*��D&�F�ʩt���E�@ ;�?��OIM�Uz��Q;wjK�����DSqm�<MP��>��y�k����f���K���Ʀm[�by��*�6�87�4F��ъi���i.���[nA^A>z�x��1����S{�,r��9C�Zk>D���{_��迈��>��]X~c��L�!��h,�����k_�
x�{d��K���^S�Rf�YB�zv�,����	�:j�TzN�k�+-��L�oIz�U��XrK���8'��"��@)9�qF�-��$�m���5�q7VI0��g�ږ��o�1d�&�� e� ;��09a�{�Ȕ�bR�1���d��2ja�-$X�&<�^����Z@�5�j�ʀ�Sk饌��qۄ	���`�Y�p ���>A�Qq㴽�}fpE�ɲ��l�j�]�ei&���d����ø��d�M�L|r��<k�NV�F�G062fK4��0��uvu!E��:�3���|�c)�D�2|M]�� �������a��EhY������C�V�W{<}�{��ٳg�l+i�TR�
�Cd�Ř͘��C�O�Z[/�ay#�(`߶ x��0�:j'��8�>�KJ[��p����M��oۼ������裏��G~�l8���x�-�_��,i�i�����r�<=	�+*+�2���G %�#����:��0��@'�ښ0�ۆ�����˜�b&6����&�C��#;
���P�L�'�M��/����L���I����s�E��k��x�'nJucr��~�C0��0$�򷉩_�jpM�,6�#�j�\��2�Cpf�!�����~ '���g��@ƬM(�2Jl�ah��Ȟ��e�W���3��?�k|�C����_�G�a��GaQ}�Y��_�O|�#��z��T�4���� �)D�נ����f���3�i;+*+�ꔀNh��Ѐ���`G��A(/U���������X
H��[���,/g
��d����*ub2�'�/�Qm���F�M��l�Ƿ�ܒ�O��K�o�"��05C=Kv��'��0��}HEG��� �̡�*�5E(	g��bj}E
s�`����|#=���	:b�R���Y6Y{K�F����F��hm @�7݆�Hݸ�-�D^ސ�^fEf�y.0��K�N�]`�0�9��5(9'�O`�y��Dr���n�����hA���������p��J� �+O1�Gc�+WobR�8z����o��'�S��ȐK&**��ҏN�玣o ����d�%�L2T�O��W�tk���E�5���QI?�]���k�@�G���k�TaI1������a�Aۦ��'� ԫ�\��u4 eQ�E}�����F��@v�ڵ�����U��n�:���M��w�ݒ[r�����i|O�*j,jp)-=$��M�0��Ep�Gi�;6��+_�w�r5�l]���u�1�fMa��Z�ٶ˪K�PG	F�d����e ��m�� -��)���f�4r�;01~I ��ȇ�T j�_R��)���5f����E~��ܠ��!�� ����c����-�o�hO3�ZOc��,;�&�UV�]�y<���ch=}�:�Yy�l%A���'19Fv��3�P[����5��K(��z�A(TȂ�ANn	��N�*�QRV��l�)�;6��a5�!�)�j^�x���x�V'\������{��ZE�Hq^��ˬ_oWr�A��T��	����X��_��ԕZǦ�l��b2a鞽{L�KJp����x	H��Fg�M�5�^�fg�I)�QJ��j��m7��]�]��o؅ͫjP�g� �a$F��r�:�G��;7�Cya.f�H0��d��T�4ɰg+J{k�֘�X :'>ſj�b�b����k2�cW|Fc�2�"�;@���.Q]�b�C�1�݌�X/|3�gO��ЇU�E�*�m}-vlj���ز�k�PW����8A���7=ˬ�����r�ǿ�y�*�)VW�*���)�����z �@Z���|Dع`�@�b���b�����e{;�`��x�]���];�B�%Hv������@�K�9U*^2,���n4�U_��
��t=M���&�d-JE/wR@��.���'N�ą\���h��3M5J��y�]rK�?�3F�!8)h�Q��H잡)E���R�|�ո��k�����$;/���Q����HP}�+o��;���zZ����d���� �O6:I�q�8 ʋQʼ�&4�5/S��S��51��nO��&@&�8qUKN{ +sٙ��<b�d�Z��q�ڛ��By^66.��Uk�iy9V�cEM!j�rPY����lԔQK��� ����[_'���;q��[$?wl?��a[� r󂈓���bp��G����$Y������0�N�����yؾ{+

�H����ڵ��s�v�����+++��7��_�mM"�ʲ���؀p^�X�ta��J�-�6����g촯�щˇ��[H*��I�^��X�إ�9�֩B����9+ˌak|t�&��0>6f�Bv��ݖܒ�O�HՖԐ4q0Eƨ�.S+/+��M�k*���Gq��QL�����T�p͎M���7�o}~��o�+�ݍ�`Oc(��EyI19��n������q�aKW"�iI;cE�?>o�Iok���QH<y�p��S 2�@��;A&<�$�3>ޏ��	T���mm=�!0^����9�ψ!>ҁ��hm:�|>��sG�q�;^<��� 6��e�v��;o��o��5"�KOkΟ9��#�d$�̒}FO�8�L�ٓӓ��� ��E$����������uue|�������%��=���hm�&�!2�\���"Ӻukl�W�Ã���E�M7\�[n��:�a>o���S��r�>{R����{����d�Yi��,����=�4���dvO+��nm�?�Kn��gr�I�]�O�𱵣Y�3�mc�+�*�*�1>܏��$�h���֍�K1<ԏ�s�؀{P��o ��!;-/ɳ�&���f0Xk�Sdh-��q��d�T[ �V�@R�Wj��xsN3�^/��l�dZb��,��i�fc�K�bz��3`c�7_�7�ن+���al���g���fV����/�y���3Ysr���x����~ݭ�i�r|�=���z��c���#`�;v �Ȁ�KIY1�I�V�Q]P
�LsqY)���d��ef�N�����4����f��J���������6�����q��Ё�T�n�/�cx��Y����Ų�\�c7�*�l�3S�IЕ�CyۄP�QS�I?�+�e �,�&�]O$(AX����FJc���=����O���?��\�?��\��x^U+���-����p~Rgo2������ g����b�H����hi�1� �\my>v��CY(���gqp�s����P]]i�R+|b�)[�9J1S3�Z9TX��p(������u�j����׏L��wg��U(�g���C�A�u6#���[�y9l�d�n[�L|����9���u�M�a�Eg5�'� v��H���Xo�d�U�~l^M�}#�*�̺����8q���*kj�}�n\s��ؽ�j\}�uعk/6m�f[�X��ڵ�]gGZ�/"Gq~k�P]V��P�6���E�y�b�lm�����A��f�;��|�;?@ղ5��+f�30�?���!d���eIt�E	��x��p�t.���౳��"�
���N��g��/}���M ���ξ��	�h?�~�8�G��ʩC[�4����l��@n�i2�l<��0CL_+�L/W�Q:���!L���7~��P��G|r�,�Gf܅���x��D]k��Z6+��x5������V����e��˞�_�<껦��e<�c�yn�@�y'O�3��E�^|���4`��>.�U�/qE��9��+yG\Y)�Y���u�o$�=^�uM&��{�m@��8�wq��V<5j�bũL3�FMt\�u۞�?���zq��w�G��;�F鞳N���pyRڬCf����Ek��"�NT(���,�9�o�6���~>W�z_66$-I�D���B�4k~�V�)z=gq�k^C�#�c��RC��[V�ǅ%gFK&�����������bY�mX�����軀3g�Z���QUY���8�d�����Ҍ�L�MY�J�F�)UZ�{p��y�f�bٚ�����7�R%��@v���%�S�B��XO�{Eq|�3Gi!+r:�l��������sg�y�m��!� �$h�1-�d��yӶ����F��\t��Ub���X�P����?p�&KB�06��vZ�j���l��>(��
ɩ��Kl���Gss3�;��/�6 �k���(e��;|��bꛜ:q��ַ�s�
�5~��E��}��U[������J�(���=]�I�oU>46`gTUSc�f��z1:8hz�����7�����#˨H ��{���Z'/��p��˫�PRQ���^�Ӹ���[�d�Y�2	�e��i!p����'bg����r��/����F|泟������c����L N�α��k
^�t��;W�t$*�b'<p|��j.�����gl�e��н���ߕ3P��p�
Θ����NIS�te�F�RJ��:�yp�5utjG���k��j��*ű躜��Jo�R�L`��U�kxF��ow��ŞH�<��2�1��u��堏g*���:�6M�E8��(;���}��7����7S��e3�rb��������:=g�fi`�L�~[�rȣ�Hm@������:o��n�X�n���R�1ґ�Y2R2��2� �/�Ʀu+Q���8���+޳g7��7`��6J���$C	���h{��-�tc���AT��fE���,'� }�C�%S&�����@�� "��koF8{o����ef�H֌xx?�:PZ��ߚ���W%zKɀyd��\O����C}U	�ڴu��8v�0�y�I3:�e�V�s�x�+_��6R�-7V,c�ZPi�CG�b�uM���-[fYZZj��5�b�@)��7.g>BZB96FF>�J�Æ�ې�8�ů}=�è]���R�/Gye�)�k�(7���dq)�<f�X�,�Ҋj�U$�,()��U���L1|��]����
&��S�f�d��P���+,�U��֖�G��5Yu��l�m�}x��߈��\v$q�a;�~�k_�ͷ܄�+W����ybL��T	Yo�1L~?z��Z��SҐ��3�
��m[9{^b�L51f�>�TYfwNc�Ro�q-.����{�ұ�ދ��/��+y��&���9��<s��r��(۷�y][������3�H��ӳ/>ט�����:w@�?Zq7��e���������t�Yz�s�[G����:��g����e�������f\\��0��4�|�(F��yn�_��]�:������8D:d6S�
kKs흖�JZ;)�x�$[�&�KJ+a;���Am]�r��M�s��3 �$g��ك��>�[�뫱�����Bt���������k+�&9�lGQ��t�e����ؚ��N��/,Fw� N�9�paec�2�i���%�� �}�m���@�t���:���" mm@�4E�3�F�S����xvFkՓlCq���u�j�����8��A��q�]��]��� ���l�S�+�*ˋ�띜 `��t)�Z$���'C�c�V�Ykb�,��.�����3��#���#�Qհ�@Yb*gڶzrb�*��-+�@!A2
#�7 � �&�U	s���/*����=��h<iR�7������l}��6�cMR������*�
�����Kc#�Y¼��w��o��Q�o��m���s�wpՎ�X�kͨ�4�xOۓ�� ����i/���c��[2x�	���M�����鉫��*��@��g���轸�H޹��X��E~>L��Ş�b��J������,>�� � ��-^=w���|��s�c���O�����.�(Mp)�~�T�0��"�:* �y&����<���Kk���8􂋂��}_��s�_�S��w���o�>�&�[���w��t\ٳ���	��3���+�	��Z�Uϔnz�V:��0AT�I˱����B�uy�s{61��k��F`auc-V�Ub66����(.)6�뎎Dcq�1�k���a��aeP�
h��hIYB��S��G=�L�%Sμ|��yz��' % �]@Iȏ7HeHĀ��^@��C��@�`�3쑭ѱ�H�';s��|�2E�ƚ2����t�������7����+*X`c�
܉R^��ԩ@]et���b�Z�)�^y��#]hifAl�V�[A6:�����
ʪ�k0�1�Y�D�̜�ze�'���NlP��!��Z���A0�Q��'0I�/�����\	��c��%�)���d�ϲ«A0,���*)IB-��c�scZ�T���.��1��}��ͯggT�xȢX������1x)�'�13��J%��Vv�6��T�V1����q�D^�U|��]�5��~��<}�[8Ծ�ߝK��t��s�펞w����M���}:��xWo�py�l0q�F�뼀��8�q����ʊ�]s�y��N;�c�]6%{R�!����Ku$�R����9�T`�O��<1 ��w�57!of�vO+D���<��[GaG�]�4*E:�o`=����"�������d�i�0�b��e�j�Uă�X�~�m�|}�
,_N����xV���vC$4�h�F������X�4;6N��d�&�rȲ�:��Hz�:%s�v�t="_c@A��~����i0V�19Y]�D�l�"�qGd
PZVJ�\j����W��8ډR�ɹt�����C)	�&��e,E3�!�,j+����쩣8z�y�Xހ{�;w�0j�� ,#-bG�t�W,�KY=����ի�IT�S9��\}�ո�կD}m.^8K"�0���1M�S��RYS�i�#�7M�S�(s|R�O�ž�粌��yp)����X���I9N&�Yx��'���K�,_��/�'ke���~3�"p�w �#�8}&���&x�Y�[�A�M���;��B��a�"i;i�ʇ^8�֖v֗�=����R�+�`��*K��<��\�5�!�U1�K���#���vº:��t�k��A�WY�8C Y�m�0ӡ1��G�sϳ����;W�./�+�t���e��M�ܸ�ۋ[ �/Cz��5�o,fŏ+�
y�����U��^�\�%�uzZ�v���ͼ2Ko작���ی�@�ϨM�*8;Oɞ�R�"Q@�:���4-�j'�mXL��"��4)�"^��G&���o�,�g*����+zI����T�fݵ�9���2�R�Ӑ��Nee5*I�t^^Qi�l����%���v��-����D���o|O?w���q��M�~�zL���o~�l�����X[1��\F�� 7� kr��M=�̇@*X�ae�GEu=j��'��/���p��w`h"����I��8�,�0�M��'�ƺ|�S�H ��͘A��2E�����x���t�-������M�5;
���v ';���JT�cl�(җ�-oz���K�8�a��Jm��� ���
�QcE�2h�����D4���?�G{vFf m�}8{�3�Aԯڀ`a9�~�Mo�'CՓ�� �]��9�k�&uH>VD�k����2���Yy�򩒨�;e~�eVuN
CU�գ�ҾޙgA���1	�姢�)/�@��=�����qu%4�,��o����'���c�j+z�����1R3�v
[��s�u��[�ߞ����Vx]rO�j�
�+s���g������F�;�񥜤�KC���أ��1͗��4蛺�<=֔.�+���fi�;7�]=o ��t.��Uf����6Ydo�<��[l91�4�҉��Q��ԕ6�圢@KsG˛c���z���N؟D^a��%���,-��oy�Y���yŤ����6�2�<\�]�+�Nɤ#�����m~����=�RNT��8}#�ig@:2|�+�㉧�k�w�Z��Ό��/�+�Aw�u͐Ah�(��2�l4+���a����rd->$�q�}EZ�;�/.ǃ�>�O|�KX�yF�)��)R�	���j#�p �?� �4V�˟�{3�G��F=�����Q<��4�\{+f�R�>��5����o�5eA�V�cv*���N�����{7��f/{�0�c�ӽ�zL�|�!�T$���s^E�ѫܞ3�)��>4:B }G��D0W:�Ex����Ё���)� T����02�r���+�d��̦�n��b˫�YC`哳ޑ��ҡq%G�9���ؔ*� S�BM̓�ِ��I�Pñ/�� y�{:JF_���f�~�Y|��'���ߌ��?}���g𖷼�^��ld�$QC6&�.S�Wv�|��d3�<
ؽs1sy��t*]|޻���9�.���.X��z��*nH����+9��B]��V��F�b7��+8�+�r6.J�+u��Xʙg7�㾧�a�}?���9��l������ �Lč9jG������SZ��I����),��꜋��2����=$�ftG����w��r(m%#S՞_�3������&�(ĕ�c�2��:l�%�tq�/��Ȋ��1)S|oD>������A�r�����<�T΀�������=
��RlYӀ;o�Uys����(�G�p۫^M�[���(�kA��4sdԘ�_b&���HE�UEe�/�q��9<���`��t9%�$��.h+LE�p �>�-�b�F����0��,�RD(Q����5�9p�v]��P>���l�s�QfG��� �Eh:}��=w݁[o���̪
@ $�̂�"�;{���??a?e&������ʵ�q��E��Г�+�!�V"�_´ف�a�$��в�	���� ,_�hV��5��(.�y��zt>�����c���~�t��=�cg.�L��@V
��l[N�u�$��+X��؀T��!=�ǟx�b\̶c��#�5-3QH���o Η,o��,�r��wT�)��t>U�T6���:��W0�d�L����`5a�S�>��������%b�\΀�i�LZʔ.�I��a+ŭNA�����9���o�Ӎ�<x�;�9��[�Η=�w�����^��w>���7�sCf�Z+b�_VW���;��'�66�U8*#��3:�(gmbFi�p������^1� A������e$0��������E��-O����t��X�j���#�`�̴[�X7�7�P�-"-ʻ.\�)�/�ԡ2\�����H��s���ð+�N/}�\nH�|��x��I�ɢ֯���7����0��gq��l۾k֬�I�Y��A2�` ��D�̈́��s��V���	��c1�k��^�?��9S��jl�!��!2G����^u�N�͟�.���)
HG���~�/����k�����#&�n*����sX���;��yuՕx�;�A*�>�S��
���7Й��?�31�~*�ĳ����gQ�l%�{G���?���,J�J�J�1�(��De�)�*],[��>��v���q��l�����[���U�s�!��w��f!ח��S�̰�~�!"(N���N�`�ݽh�� hE�
�j0�������@�^lB#�u������˿�a8:C2 k8뒕�6;�ʣ�'��,�
�W���4������u �i�s�p,	����;(�4�g�*O �X� L�JeKǂ{��ZG���
Ae��
S��X�2������B���r@��י�{:�\	��O��sӹsh�p�l4���2�v�+�~�j�c&����Ԑ�&�Ub��۠1Q%Yq�3,o�]ƽ5� ���х��"��gێK�D��~��G�m�{�����7��mC25�:��ty*�x~�s��ӻ����˥��΀t |����سG��
���
��Z�m++0�sO<����m[��������6!aK���1�*�@+FQu"���x݃4w�������(�N����Z�l�=_@��7��w�o>�{(�c/HQs6#�q����ƽ7"��pjVKM��&�R�GC�߀T��_8x�~�m���m��Y%B��i���IWT��O��L���֎g�D�/��?�<�=x��ס��������S�f�eoIt56e�c�r)Q�O��j�K���swTcV��.,r|Ե1&:�F���R�@!;�p`�d��-����_Ų�|d��,��{�Kƨ��T�deK��tYζ*&.�)7v��2N)�r�å�.$���pt/]F��8tcOi�9x�MyRX��06c�.aB��wI,Ŀع4:��D'Ƨ4ȹ��������f�]����^�I1}.���L*��8�Z������o}�jk��7އիV�S�BBf-��) 5�T|#�q��ZY�k�:#�R�����ZZ������r���k�e�U8��7EEC�������˪�0�ۍ�r�y��Xr�9���[�~Jǲ����Q~g�OZ�}��-]�Y`dS%��UL#1�?ߌ�D��%Ņ�	d���#� s.{%�-?Kbph��#���X����	"AS W�׊m��/E�2��auC5n��Z�Mx�lb��t.|�Y�è�o�p�S�I�@��=���T����O��r��B�a	�b������l�X�����ɡ84�0���[;��	�w�Pk����gP#�l�5����&�x����[�~˥����<��m��l�G�c`��
#���%Ӕ����<^���PYN���2g!�j��[6��O�M�j�L�E�~����c辞�^a%5�+y�p���|���G��}�gj�Az�J�D��&�+�Kq�x�y���`���<�:��`�q����A���<���w�rF0DOP�׬��b��[ȡ��A��{_�KEΖF�rLMP��yO�[�'�|(W�k�G>���3<���^�:W8J�&��0E����cժ��"+�j�V\s�^�J��f ��R���J�����̶���l;��I�R�2h� ����f�W��Z2ѽ�\��7���چ|�|n�����EYi9��.[�662n��<���럎��V�����Ïr֪�.!��X�E�m�����[1�m��mF��(�?x��B��D�#(��k,������Ӈ��������h�=�"��e�C*6A>o���E	v���� �ȩ������5V# �o��Cؚ$��)�^�ZV �ZJ\v��f�=��<�r-���:6T�����V۾O�e���
�ܠ|��T��Y��:��X�v	[��ze�d^r����]��1,��[����2[[�c�%�!_�K*فe�b{��֢�1G���C�?�d$s�Y��Y�e�C��8����N>�~0�>z�r�<�y	?��sy�%de��*���t�y݋�y��un��z^y��Oe�1���U�!$iS�f�u1���t_ǅ�3v]G��c�~��s>zSL�=�c��=���䣥e�{�s������z�^�,:��'��9��'�F5)���e�	M�U�5����J��o #��&UhHN�6�Ί&*�\��M��ئdc��@[���w�����Z�Ғ2� Pk!JI�f��]�+*eU�C|j��J��7#�R���ںW�]�fm�����)�e.�D��ti ��)>��
c��3�ą�n���j�g��7`+u*9CQ���ۇ�c|r�tD�����хN����8�}��e�op�]�l���l��R
�
!6>��Tt8: X�ب]i����M��ژ�?�K6�թeaŊU(d�ja0�s&�:��ʈ�,ƽ8���-�|EY)r�\|,a�M��T!){�S��I�eR�A���l�����ܹ%���[���Ϙ�RY.�P�*=�kK%����k���z��/T�@���^D{��m�7'��y��7��"�af=L=��td+k���y��k?��K<������\�^f����g�{�:;*MtJkd�k���3���U��ǡ��Ͻ����gto���a���y��Ȍ='	H��"/����m��|N7�=�
+���[�[��0�y>ł �H��~�^z�)��(�xIGg7���04<������.�/;00d;ö�������n_.>���뎽}�2��적oiYJJ�Ȱ���z�ٸ�IJ_%����Ξ'��d��.֬  6mIDAT�jbI���)?���nq�����Ό����������Pt�J!2ޏpf�lZ����)�t77�̩�14ЊI�ճ���=��I���+�I����4��������ٌ	t������P�=ڋB><���������.�r3	�	�������wx����t��EM�*G0;>���غ��� ��'N൯yv���>0k�*��V�O,ؚ�!H�p`��:��Uk���?��~�;���:|�_����Vmى��FD�I7�D67;K��o���M"���.V@˂K��u,t���ʗwo�����zם�Xo�ż��5�D��l�7��S/�04��vm��:�S��܆��"�iWWMZ�qR~��2`���X��ا;(K��g����e��y�C�q������3·���{�hcr��֡*.=��)��x��(��M罸�����S���s9/~���Q=�8���{zV��t,<��J�{��[�\-���ր�Ú�w$)J�@���@&�G��c��s��7�������m����'l�P���V\:�
O9�&��Љ_�7_jJ�/�>@���bIY96l����!>��m�&�Y:4��r��ş��?b�-w�w&�x�A��{����@��<���_j�Ye�j���K��Ӹ�=���ƀ�����Ԇ���H�)��q�E�O�g��kh@]I	?������g�3�?��D6�ފmW�2�ޡq9y�]�H��,@F0�	-�$�¹ց	Ĳ����H-ҫ�W���ʠ%�����[<��$�^�
�1PN�F��all�µ;�c��mU|�}�a׎���G��t]\��%@��؛�NaHY��?p��������7���ħ�f�.T7�"�j���4ȼP|3
�@҉d`v�nlr�a����b��Y!���W��ݢs��"1��l�z�@oF3���8`GUZ�Cg�Q�%"�x(9h�jRZ,/XѐKʖN���c=d�
S?9cߗ$�R��˄�H�0] �����D��J|U�zJ�d�I�.�K��G�@I�J�xI�G�����eC�A�W��};��eiH�/vt<
��忦�9ޗ(�0>�N��$�2�Q�E�{�����+m�_��:�})ݛ���`@�Y2�݇����I��o�]��}��h�4)k^Ӿ^JI0G�A47���Ɲ�,y_+'&"��_��t�@Z�ƕ+M���j8AL��������{��}�5��_�2�۽�~�[QU���9�(�hX��J��.,*����ǅ��΀t8
��O�]DQ�Jd�M�0��!a!�]�P\(aA�����u�$�8q�4�>��h5���ؔs�F���7@*?�2T_0�	g�T+�.��(�i�0��g~�-�����>�{lV&�����~�@��sǱ��$����PF�bCش���\����hkmý�ދ����0��*�N݇r���HƐ����B2dÕ�]P�e����o܏�>��W���2$�3X������<�dɒ�ъ��W;�=
�M5�t#Ӄ���p����N�SR�^ڹ�J�"�K�I��*ʋl�X,2j[�H]H��
b l�~������r�k���қ>Οغ�zJ�f���y����X��%�������̮��\�,Ӧ�9�>�r�Q�˧�p��ya�={ܜ~�$����c�uI�eem���L��Ιj˻ν�-^s����|���s^�:ڳ�����ʀ�+Af*�vAmY>���7���FgK:;�	���W����h���������GZUUigZb*cDꀥ�|�z��v�����Gag�]��>�%��W���/��ʺj�QW�Η�3Vjgg�X�c���������OΞE��� ��X�'9�T�?6��I6"� VM0i�5��g	��Y�D�l�:���j���*����`���ַ[e���s��Y��f���ۮ�
��R6jig�b<������Ǟ9�7ކ�@�,��J��Cز�[V�`r��#�x͝waŊ5�F� )��4�N�}.5J��HU��j'$fj8u����ǒS��W���-�(��G���=w��I�"���Xl�@j9i �Ƣ"ZhL����K�Q���8�5V{E�2��e������](>U_�|�4%�D�No��Sͥ�Ҧ�h-~���+-,�t��=�������˹�0^ӿu��)���E�c:|/����L�������=�������xG����'(mx��T߭d�tML��S����⓮�����X��3A�:0��SNCj_6/M��eN���2I8�t�+p�-�!�9���nD��%���eX�v?�Lb�sϡ���P�����ta�عs����aJw]}=�l�dﳰ̫�i�I���G�<<���r��u��2�;�>4T��V�>��}	+mUZ��*@��.��8�����g�m�aF#�Ɛ�d�2����<��#������͏1E��k2�Ĕ�E>�c�E��J��bZf�k�&�g3L,�>��>2h�'#�����?�K�N1��Z�0M������H���OU�b���>��H�1�o��ܷK{�IW����mf��J_�΄�[6%r��h�A7�$s�Ѻ4���ӹy/��w�oc9J�����G:k��������ŋ^��=���Σ�������޵����HG=#�8o$C ���-^=k�(M����x-�t|i����:�N���&F�t���{���������EG-(1����Ic�:j�T*C�w�CR�r^�}�HG0~��#��k<Y��t��ƊH����+@Qq)�**Q^Y�\������>�dG+��^�I���R[�"�)')d�}�I	��<rhp���7C�cl�ZАk*X!��Gl�v�`�+(�o��*S��ux$sU���+qdpS��p/r��VV9B��W�Ր
����/����G>�Qv~O��kp~~P~}RtVdY���OJg�]뿍�H�b�"b��ΫI����B�����2P_�k���pTyy��ʭq���X����|�t��[������DO�(ʪ��P�<�HƄ��1T����"}$���&m�^�	�ҍ5�`N-5��y�jRf��8ɓ^V�Cǎ�U�������Q�1���)Vŝ��.].$�� X41}��e�؇+_�_�� �Wpz^Q��=� ͅ ���`z �V������EvL��-]4�K��k h���{��|�]�������p� ��2,>���.y���K���?��������r 0e�}v�q�:t��!st>iCZ�*=K���=��-EU砣��a>�����LY�轅��O�S�[�^d�x�i`��4h�%%���f�Ql߸�a���G��s��sfS��TO5#?6>��"�K�vg(+/�*�I<�^[]Sm@aՆ�hɨZ��H�Z���Oa6�����f�زaj�
旌,����n����i������{G[��sS/dF�c���7�����)F���s�:�7	85P�E����ᇓʏ����^�/K5��n|�91V;I[)�������t��
�5���ɴ�1M��c �P'�e��>��!�J�u�*39Vr�����c�,ͦ����X���<����޻gN�'f�K����O��l��� �▷�q��0]���]#(9`bc�w�ֳ��w��|���Sv�v�/hPy��О���I�R�X����ӓ ���x��w��?R������p��^�Y�v]��<J*s���E0�	�(�΃�җ~���g֬�G7����	P��ҳ�.�¹��_鱴�Ӟ.�ij�[�P��Z0碞b��M�7�ay#�1���cȥ�YS[kL������f�|Ŋ( ���겭v�***����,�{N�Q� dR�1Ɂ��:��s�Z�K�_hg@*}�9�D��R@�òX���!$5���s�G��!�R�a��YY`s��9S�C"��(�3*5��4�O]|f�Y���"E{��=�[;�S/�f=c�azLdɲJ,�W���̰��?�a5�1�"ښX�H)}Mft����?5�.���;5��iAB��(	��U���Y�u�Y:��z���Gu)��rj�O��^������������C���Νw)�W����޽{/v�IG�h}?�/��Y��x3.c�<j��<���h���u������^�ӕ��٘;_�<�8���b�㵴W<j��1�xC<*uJ�E�o�{�n��_�����I�{ﹲ�gz����QD@���3���'vLL��N����PZ���UIr�N�����mۊ{���xV�^�R�U�� �;�1��1���c�8u��=j X]]�4�����hiif[�6c�ʫ���c�T�����:�Q{d���->�Es��N��団�09��`/&{;�n�8�H�y���P�y�^�h_Fz�1�ք����t��g1�y��[0�׆q���V>ۊH_;��݈�� >ҋ�h�c}<�עC]�i;���Rw��8J��V�=U��6����D�=Aj��η1�A��C�%ZkL��})Ujwԍ���Cd|l�d�QLƢA?ӣ�`c�E�T��E���s<��ϳS����	(�J`��K:O��+����<.8����|H�c/��5y�A̓�=/��`X������(��s=�8\��.���+���oƂw��۳��t�.y��K�����Jܖ�Op����U���K�����T�Ф�I,�� Od�4o�<��;�����h,��LCR����|k��Ȉ�B����l�y���NgϞÙ�g�S$Ea��z��04<d��j�R��51iݗ��t�0}�����G�>~:������/�c� ���2�1� F����DO��Ng��t_�pW:Ρ�����d`� 0N��#1�K��Fd���-�.�K`�yo�i�������3�k>�ދ�	�'������(/�5�R�t��%��$��4V���G�`"6�s?�K+ػ��4�#�����w_l��P6��Ӡg�R�����U\�X�1b����ڕ��K��E�����{��ڕ���|Lo�K_WZ��?�y�"o߁�=K�1,�p𚁩DY�����=�����.�(�t��TuL�6ϴ��{i�|XX<��wa���5�K��r�(_����O�K9�gL�1Y�ߕ�{.�� I�� Q�w�ty�&Z�<S�������k\׌��Lh��l[ط�#�irI�.���,:i�w�i����-�m����5LUX\�(�-���$��Wm�L�Y����c��eƲ�A�ȿ��Q��2tf��}t
�����ڎ��z3f���D��@c�R��f!�&�I�B����4�17�y}H9�k��UW�N�ߔ�Ĉ�r(�%qӵ��w�U���Z�����9��7���	��j�21�t���l|W����5՘�@o�lX�k��A�-�c$��4.�R��t�������.�V7Y(*�qV�c�ϡkhMm�x��$f2�#���d��e��JMGb��5��1*:F��<�a�y�[ɣ��=�kL���e���S>�զ�	?��i�A��{�����os��g�4.�W,m�>��ml��Ĝ,-���N	�	.q�4x1[��k���U�t|�rn��N����L8��=�-�>ū�p�ö������pދۮ�E������=�~����¶��s�J�o/��+|��6o5�6G*ҏ����ͯ����7��������)9~=}�flD� ��{ld�f���tҌAbhp��/���u��׬Cs[�mqs�ͷ�v��<������W��>��t����w��n\}�j�\���VY(�^F��-C�A��vG��O���^{�]X���h�,i��c�"��q�96�Y�� �T��	�8��Ǌ�^�����j���BPY�L�8�����sx��?�Mcٺ-���	���=��WS�eYi6vol@~nz�ڑ��k�ƚU�L{`>��Z{���Ng���Ջ����"��8]�/��FWE;~�	��g�A�8߂}�C ���r�� ��TKC5k�u��Vp.<�8�t�\e�.]�)]����G�R�6�6Psૼ���H����4|:��Y}��)�3lE�^]ѫ^����G�ss�F���G���t%��<�󾹜��=��KBX�>�/]���(�(Y�����+�ty.�"���Ώ��+��^���놃~��R��������-w���A�>׋�ͭ�@/&ZQ^a��ɨ�d�����PZZ��`Ѐ��$E�,U��U`�b|�� ^��7�$�Dl�������$v��&���y�,�Hz�ʸ��o �_: �g��82gSd���2C^�e�����3���cޟ�c6B,��?�X�|0u$��'�d �e�Cf��lۈ����ȗ,�k�tm7�^0@6� �Hԡ(�I�y�?0�`n�i
h�M�,D��Z�78���	�_��jDb	�on�E������j����//y��.}��@�F%���Ȑtl�;��F$�DGo����t�ӟ��S�����z��"�u�����~؋�\��[$醨���aM�F��o�g<�3��������$}p���n������9/L=����<{E�8��zj�J�,�Sm�b��M��;��������1�4Ѱx�㿅�p�\�i?oᷜ�c�j�w�$A��*�E�3a����eU碱])�Ԥ���5{�D[�k�J��!�Ei��$���ǉ!r
ǶAQg��g�(�SMj��:�6��lj
"�2I�6�D���b"C=3?��-]Б��LğK�(&(��s:�����k��bO��w�W�j�>�&h2��+�'+C��݈����3�J @��fE�A�Ij��G��(�B�
��?���N2g �zB�H����Ѓ/Q�����	457���c;z�1HQIiqk�U��d�@�`�Ḇ��m}5�΍q��9_Y�~e����/�/�mx��Ӝ�8�<��F/#%V9.�]y�w�|��9��������;a�1��/����qe�8ޗ�
�����ig��F��E��{v>�i��x��t��^����;w�?/�w]��PA�Ĕ�xc>�nb�dD��`�te'&���墵uu(*."��*(Š��J��q�
466�%()�[*��Ɇp���xzu@�_Vg�0�dKS~Dg2'�&Üc�Sd�1�O��dQ�&=�� ��T��,0=;�h�}�Ӽ�$���}�C�8Ï�"���������{��&���2�!����6�{
�f���T14��J#��GS����wh�v�:We�2�0��.\@gO�ͨ�k}�	�DU]��3���{���l��A}�a�G���	�ZPJ�>3�F��h�Ӎ�W�4c|��u��o=�g<0��_��{�=B�,=ʰ��+mN$V�q�{��?���떧?�v.�t�{��~���%�{G[�1}cׁ��G��<��,,\w>�Gx�4�.��c��LKE�o���yjN�����B多�I��ȸ�?*@��|&Ύ_+�d����yZ}H��-Tr)����ڎ��������������&���PN���:E	W�r�]b�6��v�I�%q6��2�?���#�ر�5�������uj*a�ULN�y���+�����Jf�9���T+4s蜞M���9s|N�5;�w�Zb�t�����G�F~Y-���|/>�i]@��L/��T������c�l\��#���AMy)�l��|ղ��K�9�����F����3���έǥS�F����'0<9�I��3��h�D.Ӝ��Qϰ�d֏�ո�lF*\���T+4W����,>W���u'�L��S;נ�{3���K�u+	�ty��50�K_�?�~@/��?���Q�������<\	����اҡﭔZ�w�$�:������id�D��1�|^�G�-Ƌ��-��8u�.I�]y�˹	��8��'p���p��;𮷿	kVԙ�U_o/Μm��٨�����HDI��ެl�f3L�;>>jv��CA�8 `, ѩ���$���ӌ0w��n3Z�o�~��_�/l��s��~�6�j����^��
l�t��+�.��H�]�q��������/�#c4�Q�~��N����V�D.���0�,t]S�\l9�W�Q	Ɨ6�K���V���N+������D�,yj+6l%lfab���:��iX�;�a	�5�T"�ʒ|�ؼ5e�������-[��n�o��5-#�J�kWt����B��$@F��Ԅ#'Nbd2�L��#�8N\�h�<����<��O1Yz"��B�����9k4V��cQ=�u��� /���/�^���41o��IH���n��p��ҙ>������.��wGs�;I?)�~����0�N�m��gp^�p%��ol��ixy�}!%���s:�:��/��n�/.���eM�v&���3V��dmP���k��ɞ���(���s�`�:����N�W������S�d����BЗ�$뮆�f؞R�Z@3C�U^n�b|)ϓ��0]a0d3��{���!@t��C����[l�����d��3�j�*����Be>E|��H���#�H�pǚ{ Y9y��S��Roߐm�mCF�{4�#AV��|8��c��$&ӈM͂�#>=��|r������&���|܎�zw��Ï7G���C�ͦ�QU��Z�H��;s����	��d�qD|��xl�b� J��J��ؘ-��ɑa	�v�t`j�̾�K9�����J�q�6V"�������h�s�nV(����e�������Cz��\:N��W-r�-Թ�{���Qz��K���u�=��9��7��L�K��ĻoC��y�4�[^��ӿӁ�~c�Y��]��.��8�~{���e�j��{��⻜wN	��,Sr's�������K�U��K?�������Q�����ȹ��4)m�u9��{Va����m��d���B|b��
7�[������wvX?IX�eŉ�nfZ3��U��i�Z���$Η���r���9��������$d�Y������DA�2h_�Xd�uոj����u4g+�s��b�v�N_�.c��ck����Wݹ��uq||;���v��IӴJz!Zh+(UC��J<�E|'� /<��P�
���/H<T��M��b;��\|�������OBR�JH����ۺ�̚�5k����Z���;���r�זW����R5���_*EcӘ�R*K��j����f����ֻx��$_�������?������=xX�qʋ ��3��L�S���起t�.�8���bRݑ^�V䙞>�$���<ӹ��X=׼��Ǐ��O�����l���pC�n�t��yΠ9cL=	`�݉/�ǟ^��6yh.>���]���f#��2�#2��d~y�;�ס#S��Μe�udi4�O.�2�G�V�/��(�r�?�_
(�x�?Yh]��K�\�も�! ��cL�������J@�W<ݫ=AxA�*4p��Ϗ��o�, ~}YG���LE!����#u�[����z�"&L��2t�5p�G:l'C1��LU�����=2��9q2��Ix
� Ƙ��-���7VcbO=��F���������������IX���CFl����bK����v`�2�jm��ʊ�������ː���҉��O?�>�_��7�'����?~��_�ҹg�m��W���g�����bf����e�8`� =�ϱ����lH���V��FW��>2�bl_B�+��m�bT�%���	���8�+X���� �j�8�-3����T ޕn"�a�8W���B��:H%��QDp���6tO��c����̤>~t�c:7݈��zl\�SJ~��8%�:Ǯ�ӳ��h*o��B>
Fp�Mm��K�-�%��P�V���ťk[1i�<��*0J����B`�B����h]������?������n�g�[d�1���N�����@ϪX��d�|^N3ϼG�% Q/�n$��0�6� ӥ��}�=�hi��#1��9���C6�_˸�W��9�yH
�R=���(H�4_��CP}Ɗ��:�`Q�xWH~�s�e�𡮙��W ˤ+��ZJqZ�EY~�#|�2HtE���רzm��[1ۜ�eD�y�I��6����9(ٟ��NV�!_,�w@��u��I�U_5��$)�R9u㷺���rz��±�8<?����x��wc������W�Ņ��ߋg�<���z�J���#祦&��h�':�����_W����9Zj%.�.��o�h�2�=uY˴&��UF��^+K%��!#`%|������sB����:���Pz�veȉ{����y�	Ϯ*h�qR�L��ڜ���9gU�������^�+�)	Ps~)��g���/����ӗ������7�-<[�AK���My���֯�w%T���/լ��J�y*����9��� ���gyا܈��!S!(�X�n��8���'6]�8T��݀��P�8T��G���Hg�'=]@��X�*H�Ç9���i���q���n��d�O�����Ҹ� ���#a�1�p9?�)מ#*��5�P�4���2��FN��gDfՏ�3���'��@U~	���]�OG�`�-��7�%>ϝ$#G<Hw�,˽�v���ci��F\��r4g&c~����ȅ�H��x_�����N^[U<���ŉiy��ɍ������G_]]�љfl,��Sg��k/��Ǐ���d�|�K���dۆt�a��Zx�f/~�֟bU.���c1"�{2 �L;��:gY.i�'B@�2�wLLo�ʱtU�ܣ�Y�ѕ��9`o!r���TR��
5�:Z�|���/��<ط��%v*C�L�٣T�����@�7���q�����fV���v���;my�c��FD�Ce��>J�^B��*a$Z��ؐ�m�����7n���o�.|�1*�_�@/<H�c_X�GN��1d!:0��X=�)	%M*<�8�aE���:ѽ�#�Б<��;����x����:�2.̾(�l\�ϫ8�t��»4��gj�Z.J9����]�
������F�4���?"�t����s��A�Q�q >��G��l���u:Ň��L%r��0Q�@�f���2~刜�gU6uc���14�>㚄�/���ʏV�`E_6�cVXC���q����v�\�Biv���t��Y�nl����1�<��I�-ڥ�����0Ɠ�GhU֎d�Y;��gc��Q/˷���9w.^���(T�z{1iK�KeJ�����H�⍷ގϮ^�1����ї �Y�zG]*��#��(��I����T(��:G�m$ �G�9���5���'����vp�9�x�E$�����8�5ʆ0�nĻ)�[�jz2��qX]�cs2��V�D�s���8����."o+��L��$뛛�:���q+�����V�c�;����O'��@~6~A�1%�)
��|����M3|2�Yћ�7|�������.���<"��G����0�ݰ��������*W�3n��3K��G���T�
`d��ң�m�PYVyn��P��. ��2$>���'��KP=��?���$��n�[.��<_�Pf�,��HC���,d���s&�#3�B:����U�TW�A�kF�3+�il5�ձ\3հ�//)�@\���3���уK�(fDzB��n�۪�w2��zì�<�uȻ��#G�מ_���0,;���B<��;N� ڄ+s�N�%�l�r�֮\��Ξ�W�Re��AW^1��H�M�wȄn$I	�x�'Wo�_��G|p�b�n������}y�^�V�W5C�q�] �
C1w���XwM�J���E�[*���R)�TpudD bAAHK� x��eAF +]y�Щq	Ä�g�>�X�NLN�&cS�"�'bJ���+��ȨT�7u���Qw�7�t�vpP�j�y�ٖ�%!ّ�l��m�X&>O{x��MDgC��`�ۘ�w)� ��JHr��p�`����ś�T E��䛔Gt�͆�����׹��x�(���1��5��y��Bdh�:A���+F��(���3g���}~�#o�Y�P����}�z�E�cy���r�9��i�<���J��m�J���y-�A�<���!܇�G���!�i�#i�'���V��#V"�/\6?�+$U�� }��v't��o�c����ft�:P���`4��ȸ(�(�y�_�2��!F��o����|���������7��7ߌK�.ǡ�Y�;��;ۦ��%�Ӑ�cpY�yzj"z۷<��[O>�������c1'#�l����I��ȋ ���,p;��5�����Z�߆�owb���sŤ	c�|>
�R�	�*�����b�|PZf\y�(������4�*��V�J�.Or��g���ff �D�L��� �[�\W�
G	��5�����71��Ŵ�x�gyF�_IE#�LOz�Ǧ<M��n�r�[w����<t8���P�*o�-TXcA�w��֒u���H�0�LE�K�a�-#R�P�J�2X;rO�R@��e��ep"��gG��=��
�~,�������p>w�Y��S=����*���$�|����_LAa��^=�L�۠�+�������?i�y�� z�Ʋ�F�x6>*� 0f�Ƅ�	/�|��F�x����-���ĩ������q@�'N�T��"���F���	�Ax�^�C�y�u�^�%+\�� ��/�xn�Tw�c@�Qx�R�DH���X��"q
���bZy3���;�Ϭ��|��:�aȋ��9���C���/za���}�����^wY������c��_�S�����W�Vz���S�+�Fc<f���NƏ^�n�=}*gZ!n�/K
���|3!I} @���ޠ��/C�P%
y�(��/\70<T�8z�ב�9�A��ÑG8��p�y�4�
b�:��6x,�w@%S5.�폎�82�����@�����"ȴȮZZm	��9��e�Ɣ��d1^�Q8��`/�i	�H��ET? ��)OQ��A@�QX�h���_��d�M����(;��Ԟ�ۀH(E�HQ����ޠ��[�K�GJ!%Q"N��w.@��.0d؞�;��Un6 �:D%VP���b,�S���p2cW�s��Ҫ\h��r��顼ɧRe`��j8%ƬU�� ^t:leC��x~2�2$��U�{3��p�T�28�S6�J�;r��7	ʺ/9�`C��i�uE��䔢*/��^K7�n�[�L`��C*U�=��3*��M'�i��rA~𹭮~.�ܵ~l�ߊ��u5PS�����֖+ae|�O^>шRJG*�`a᫚���}�kvf*N--ʈ6cFeB& ����o%Z�����A�T��g	r��~
�IΓ�}�Y!RG��j$=�/@�0)��#��YPr�_�O�x^L��lVހ<
�	xyĕ�0��Q�8��F�;�S�F(R�	��f
D�c�һJ*Jɳ��R�W�Y�֯�|�����n��z�.0��+P�]9�3Ɠ�Qclm�t]q�*��C����~�`Li�H�+�AP��m@t�����Ѫ������^�,Fe�@� �8�G��=���`���lx��2�1�}>`�o��{4d��q/�.y� ��Ue�6�7�(��J�g8=�Q� ��0i P&y�y� ��N�^�A���A��� �	�L�h�    IEND�B`�PK   �F]Y�'���U  �U  /   images/79f1f6d5-8698-44f6-90ff-b688d5ed2669.png V@���PNG

   IHDR   d   �   b܉{   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  UMIDATx��}x���ْ�{#$����+v����z��P�]�a��{A��bGADA�@�=!���ޓ����̞�d��BPr�����Yvfμsz{ߵ�װ�6���T>���d>���G ���e4�Q��j>~���5_����67��	ai������� ����������vt�� �W2�S����|L#7a  r��0ANmG���4�	��C��Z���L6&D��J�� a����FA&�A�csP��������NN�� �Z\��i"�1�����L�����X�b�	2$�x#۟	0(����Sjx��7	A��a���]A�E�<�\���'������?���K'�5,z����_�_�)���7�Q��J�h$?7A���)�*�V����jj��YF��A|L�)���U�^6��n���G�fdQjX5Y�N���>����Q��2:.-��0Afm�MKb�#��K3�7?+�D�Sr�?�DPB�E��Qp��l69�ںF'��4Sae3�5��D����jr3���c�uTc�-�3zo��Q�"���[��S��
:*5�r��軬Z�+Iλqs��R�(L�Q��L�`ѻx����-*z�f��r�0��wٽ諭}ξ�C~dBL ��NG�顔�D��ڴ0��]�G@\�4.jlvQym�7R��ZZ����m�����x�>G���<��:�W���	j�k8M�C_7|a"~�a 5�:3e=�՗�)} �q=�<��������k��F�g?.��b���rV���j����n��e!�"�蘡Qt���th�0�����p�)uP}��8�!V�?��J��@EU-�dK5}����.���f�0�=�R��Of��Y#4��6��q���Y�G9�3�!`|��C�	G��I��_^5�L��_��U��J1�@H��h�:�����O�-�]>69��;�UD�Տc�9�	s
"B��7�w,)Л�}Qp+ssbB ]rT]06�z'���w���ڗ�q������d��FE҄�Q�]�H��QB��Z@��{�~�S�ل&Fe\�g�O-k���H���G~��%b$������z����^3T6�>nAz����a3��T�N��k��,��~�/7�EQa]0���k���|͍/���7=���*n��ul̶WDvh�E�0�"#�����c�>ة��Au�F�=���`��h;�}v
]qL�;��^��Oe�Mb��� �t~w��B�B\w�K����Ɯ���ugu(%��W&�2v�ίh��q�*|1�8f榥y)ʰ��4p8���y1���7s�B)�椬�zy��������3���O����m��G@�Y����^\yP;Ĉz�qΑ	��T� ����=!,�)��&�ElH��t���p�_�?<Rs�Y)t��q�����"& �Uc��x��2+�fZ�_�=ӟ�I�EI}M��Q�-7��0p^M(E4�	ǚ��/p���.� ���,�����g5�yT@Û�5ad���۟m�R��X�N�QQ;�æ�$�c�8��4��X
��c�O�OB\ =zq/:��h��#��n�*��������(**��;w
⛛��������)44����(==����(<<��'6�MMr������=�l��5}�Q1tׇY��՘��*ґ��>ޥ�Mf��,Sz���o{�ܗ1��i�Q9�=Bkެl�?�5ʹ�1p�g&q� �P�8����`�Y4��5�d8�I�iw�_~�&���L�g����@	��XETc܈(z��ޔ�Sm'�	����/����i���x�bZ�`UUUQEE566R`` 544�u�����'D0` ��ۗ;�0?~<���l�ev�x���h�3�d�n(���6����U�M�!�$xG�+4���>�[��~�3����f�9΁�\�BcA�0-D���U���P��7����#ɗ��.����Q�̱[���rc:��8鲓��ы�ȟ߫#b Y@,�<w�\�1c-\��JJJ<*J�b �AAAr��1�ÀĬ]��V�XA�~��H�رc��Σq��Qpp�Л0�Ja[��-��Or���
(-��s^f��qVZ�n`[�����L�u,UC�k����`�ǁ PWH� ��h�aI�Z}���}>=��)���,�l��Iڵ�C�H��h�Ѡ;�Mc]݃�[���jw?$H�ꫯ��ߦ�+WRmm-EDD���H�-//�;�k���D�������BBB�p�����?з�~KC��o��N:�$y.$�<��yl�q=�OV{�<��Ŭ��qYv�.�+�*��)����~��y�n�P�R�b��_	A��.�!���<�!���6��F�_\���\?"ӱ�0�֘<s.5�=�Ѥ	)���B^)\�C-=��C���)H���jH΃���f�0����R#�����^|�y��ęam޼����
!���N#G��� �gs�~zڰ�PZ���,�u��t.������	�G�~ggxV�=iq9�W�7�cۑ�ק�3���K��,H�	cGӰ=�����y�z��gEB`x���dH �4���������9 � ��!��p-��	��1�|Hޏ?�H���q�B H�{އ�k�:�����e��E����/.����b$��pʱH�ǂss� SY[��%7�N�ή�
h���CS�����S��ݺFJ�MeNJs�4SF��i��0�%�������.��o���P@��xp=��.>��wv�7,�E���{��iѢE��O����<D�H��E��U�u㒴���T�(Y��;��'�����B�uH���6���7h�\	"�_�Yہ�eS�b����x��C�Rr�=Qbh�P�ᴞ�t��%����Nf�w�3� ƦM���o�e˖	�a����h���'�\[�Ϫ�`3��TeFii�Ge),\.���������ϧW_}Ul�zoJ{`CG�DՕ��;vl9���LRH]7�!ze���lrH��&���|��8G@nqg3Z��|r%)H�p���kg�������6?/�f>3��� �.���ǆ��o	
��9��6?b�#�ƍ���/]=u��g �[\\,Hr*++%���
2aԨ�>� �-,(++����Jz��iԨQm�bH��F��@�U�߲9;�������7�� ����ި�soz�ƥ�bF�Н���<��)�n2�C�Ȇ�������h񹛍|�ؗO��	��,�����i�Ի�!�g���wPbH!q�N�����䩯[\��!#����x��m��%��^z��<�	b�����(p/l����pi�X�W�ciP��πc�Z���,H˶m����׿�6����4||jMM��7�n=�g�5:���2.��5�s���E	�;%v�	������pJ�K�8'SZ�C�
&���imI �Q��PV4�|Cl`=�ԭ�o�6i�9�U&���|fR���1�1�tp�7� /d�.7s�9b>���6����3����yH������믗�R���{�eD�vn:�i�f69îir:�6�qc���粆�@��	�[n2�m��k�^�&���T��/<��fI���&&Ʊ�O�cvQ]p�c�Nm~����=a3B��of�I����aG����í]�d�x8xy�����32��U3j3�Z@\p<�{p��竗��8������=��,H���/�u�V���E}�'0��C%��g�57�pڞ��˪ƀ���x�G����OtX\'�wuK�e|T���Op�tm�u�AB��'�o#� �����j�8s_{nb]Bp]8뿞��@��`.��;�"�����z�pc�x����P-xIE
����:D�kAD��ǂ0J ܋� jJ�5�PkfX &`� PI� T�|x�������'P]�I��{$mY�0�n�@L�����J�fܤ2n�<�eɀ���=]pLd�۷���36$VStF���Q���Q���j���L�m�]�N��6m��w�,�4�J ap�p� &�d1@8��yp8`�>|�q�UX@�@Jp�{��\@�G}Tra�{�n�8�̀��Pn�*&��)�qӯn��
8=�m�/Q\� 
 D���A��ȟ�+���S��1�[�S��j;%g̜#1G[xz��%;�ċ+A��P'-����b�gF��@����q:���;��k̰px��y\IB���/�Q].�C�=�Ў-��d�����D)m�VDj�C������|c.�ɯe���E���+�
u=x�l����e1���")� C;g��8����S�U�|oNwh:����J�8���{ ��5X@4����p*��;GaA=Bj`�/��BQ_���b&I:��������)>���oP�e�TE��5���{���iC�NamKA�
�끈a��Fcz�#Ж ��O>�D��*�.�i�`���kq�Z H 4� �{�2q^��
 c�a�&��+c@Ͱ0�L0�~x)i���Au���J��7z�_���(;�8D�������D8��H
�P]c�'�E������E���������������j3��8�q>�a�>�oX@��;oXZs�yi������:t�癠Kp ��c"iņ2���G/WӇ�3A:������`��v��Y�f	7��Rxq�0�p�&�=��:�os���&�<\.V' �`؁t�ă�x�8{����0TM�4p�A�1�x���)0�mV��KMy]&9\Էg0�Idc�l%^
����/�E�q�4�j��8j�[cU@��Ps ���8Dai���t<��1�!fX`���k�����t�m�y���g�� Z��F�W�ut� <�Q�`��&S��@�
E!�<8���!�z���*!�AB�k
]��r��u�R�VX ���́`g�p_G��a@���#��H�D���F��U[���@��Ȍ�v�A��� d��TāXu51���s�D�980��
oX�絑Aai�
�U��/����B����Bou���Kg�+�_R�T��/�t�RA$��Ѥ�Q=#ﲫ��$���p�zY�*_`�:<�j�e.+,�� U3�a��5kִ�!���}���o���jG�&!<ш?J��#���u����v��Psb.���2���q��,-��3,M�h�y0�C�fh��5� ,<�W�Z��0���'E�-
�QiU3�+E�H��P;E��$޴8��\�io����d�; �Ƶ��q�Z L3,mbPX@�ڟ=�BU� KEoX��&u�A�^�zy"M�mF��Qi�^Uv�/A"���&���?�F�ܚ�ut����f���Bu��q|o�����<��`��|^����Cn˃
F@ �!�ԨU	a�d��hq�uy�m�D���,�ЂH�9qʙ��5�pa@����նoX���$
כK�j34��W�½�K*Q�?��Z<�\��
+�+����>�.{Y���Ƶ�@�MZ��|��!��5�.��Z�̰`\����z 5c�i ��8Ĝ��PX $���+�z�[���2A����jt��|�������|��p���jP	�*, Mai
�#Xj3�a�������7,M�(,H�f�;V�_�+>��.����ƻ��]F�k���͟;*�btT����[��RpG%es���̍�d��)->m�ä�嚛Ҭ+8S#dp ���v�쮄�6C;E�s����M6�R��,���l0��:"�,rvm�k	bq{%�VaӀ���Q��]v5�p���+��6�\���C̭�澬=�R�5�,�T5�x6��]8�q�7���NyX,v���ߘ<�d�4�in
ÜqՈXcp�f\���j�ޚa��WX�z��zh8��R�5��gs�K��j�[���A,����no�Y[�5�p�sg��{vt-���Y��g����Ka������Ҡq������"�"��Nׁ$3HL��t�X�۟(�#p��C�������nj�DS�eWp��3,s��̩��`�K�8�A
�fx��ԉ9��s����.�d�e�5�W8O���C<߁ x�>}�Ȣ�����n��Oum��0�4�g���[IͰ4���pԧ�1���,z̘1�EE���xH�G��~���5�p��?%�(0���=�K�u����ns�>knJ�|g��nW����y��W=X沫��a�� ��XZ�Z�"�ށ���K���L�3?�Ġ�]�i�QC�c≉��0S��z����ԶRm�Q$j[�X�#Z�0�ҥnfX@��`���P �&T����r�"ARP�5����&VY=�äb��٬}�F|H���B�����A�  99Y:ȡ�4��]�UwS�����S�|G�ܫ������toX ���kv�;*�J�X�سg�v�#3��-<���6Y��/��B�2��R鞐S�3�<S��A����Z���E��p�UH����Ͱ���l����a�.e��qfX�r��V -�{����fP{h����,��還�ʲ[�nkMucRxU[㣎:J�����
��n7��;M��ZQ��:��DEFg�4Ů���,�Z������AG}t��	�ڄ9�٬�8�G��%	�����Ĵ��CS!�]v�,�Բ+�T�yH�6�A�h������b���u�Z��`��, �kw%܎`ib�#X`��/�X$G�V:�a��vi���2�DY��V� �-Q)�wg�u��7G�d.᪞��4�����fX��̰vW����c�,wk�FjzgI����SW��}'?���!K��趵tk6��6p�\{�m~jԕ��Z �C�@��4��TB��*Iai+)`i:~w�p=$\��B����`�"�q���K�kpP}Rr:\��X�,%��v���3g�i��*0��.vw�î�[u�8\��������O̰�<��g),�
ש��w��駟.s7��V�t` ��Njlv�(ᢏ�=�:'Ű1kq#XS`(a�L�"�A�>д��eW]���ZT����r0��*]�R3,�i����}Z��f ���&K���8�.��U��UNr6s�l��	�y����e͔��'��i���z������TY'���;i�C���q��J���nn%5/i3Â�0��.�ai9���Ao� 1@H�V�*��ܒ&�'��qE�/#��`���hlZ UT��գB��/u�1��c�=F�&M��T���W���U4ī4�^�&��0��̰��+~A ����H��s�p�	m솪*�1�q��+������*��D.g)���z9H�h+(���z@��?���ǜ~�,*>�[q̩v�sJ]�e�e>��|����W]uU;� ��^�C��=���YT��u���Jj�^�Ni�*#!!��=��� ����/�=�]��4uĀ3�eWݍA3����6���j�3X��0��'�ۺ	��֔q�:��YBv�H�u_G��]PK9eN
�W{�L܆���֡D��|�Ѓ�_�j��:Zvմwg%\�݀�%\s
]ai
���ӧN�*K׼�x�e��<����M�,=��l�1�D1��m}%�?"���+�MVS�VI:4�`)�ɓ'�FcZ*�}��Gm���Z��:쀶�`@B�\��6��<x�8�rH�X� �̩���¢"��]2�]_��R���B�dl_j,,��`{�� r��x)H�م�K"M��g����������,_ޗ��6����T�u�]'N�wZD��dtFQ����?�f�Xo4�uat� <����hG��,V[�(r�{�2�cQ̆
n�.&L����O�s���n@j3Tei���,H�w	L�IL��AH��竚��]����&�I[r��d?O���sԷ�����qqTR���$���`h$�k�.AT�v~��H�{�'�}�y��7o�����V�*\5�dM��y��- �B�	�#�86���������ɒ�z�c3
d5�Ŷ��
c������3~ͥ?�j�s� �wj7:�*@�Ð�U��Q�,�od��ٲ�oݺu��LW3Y���^�v�@Zt3؈c�=�N<�D٥T�|ޕ?]���;�ax[D%Ma���u�����0�A�=wAa-�ZVF��N��b
鴵S�����F��������\s�������0[�l��{a��e��a!9�V��K�H=z�h�,�{>�
��׾�N�Y��u��3��������5���?"����7�����NF\X�{}��"aW�� -e�S.Z�R��8��S=�F��3��s4��m4T%��B;�̼'b`���E��hz��?DK쏱��m���k�_�쑽� /��⽛��]� �k� 5c��5��b��Mn�-:�{4h՜�v�h����e�4�?������?ҁ��$��d���t�!c�ΑG�����\��n n��h����)���v4��@M��䠯�P8uuh
�%����9$�B隣_	[R_�DS��@�\;�/ZHCz�e1a�M(at��zT���6q�r�ΆJ��� ���!���7����b��Z>��05������ؿBX&m�_��̃�����i�ֵ4 #�{Y�TÏ��w�F��fOH=,��ɜh�W"�@ANA1:���&�Vo,#K�����N�1�|���}�p`S(g�.J��n-��Cm�y�t�kj'|1ξ؍��BJJI��;��ܗ[��/10��@u9�t�������d�UD)I	]^��y�Ų[��?�kWA!�Cb��L�>��{��Y����ϱ�eL�wL�.X����҅Ex�d��*�&k8�N�n�������0��� �'�6���ϯ�7oCs_FM�y���L�����@�@�eNn>5�EӠA��ǗQN^���_5�R�`�?_�YLWL_Ao�|0-X���7�Р>)d��wy��_1�R��D���)8:����O�=��6dU������	��,Z]B�?��޽mm�����Ө~��	��P�TSUI붗P����/4�&<��v��ˉ��DY�UI'߷�^�8�F<��/ZJ*�'{`ZZT*v�R^���8�(Z��H���.w��B��� 0��Mt�#��s�ѥ�K󗬣��iX�H���f���I��X�l���ژ[I1ɽ��c�ӳ_eћ�eI}�b�kxG�o%r^����7�O+�ˆPȀt�-a;�h@O�ߋ�����RiAR����UPK@>��.q�/��۫$%�7y֞�C^�#�U�+�Va�ӓ�?uUTU��U( +�z'QBl$��`�+��1������J�i{qQP�u$�lA��g[�y�=���� :��~�N�/�g¤��GL.���ٴ*3�bwɲ��$�Dr,�<���ם%f��$"��A�*o��ՎK�A��N��6z������Ԃ_��TЁ� �W�F���>k���9�x��T:l� *)��m9��fS1�e��`��Q`�]��٬�jѭ-�z�����7SU��j����B(&6���H��PZ����|���.��!����
�8��!`�=p��c��L����Ó�A}��梪�z*������/��%�NI":Erl6��*��J"�(4$��]�aG5��c>����JK�C6�J=u4�At�ĸk�e����ɜ�l�4&P�a�7%�z��Rb�?��e��o����3�ŕ��a[m��壚r��C�Q7#�yt;������[� �[v�Ж�j�l?���{�w���z���J��\b��e ZN=O��'���Kǿ��e����C�l߲���⃟���Q.��[b�����{��0ͫ�D���7�mG��^X':_T�^��0J���������(�%-kW-mɯ�#��v��I05[c?^��!���+�^��L@�����*�����l<w@Zm�UG��FR\D��m_�SE;���nEy?~˧�B�!~�ǆ2���T�0&��xk������D��7C��iCV�q/���[�\̅���]�������#S貧W\
3�����;�������;"�wq�c�h3�\�g�L�]���`?
b��/�^�a;=�lK]�n�ͯ���_x������tۛk�Y~��K�����33hқ�h-�G�"����;��{h�������S��Άx��:��#��O9TZ�L5;�IǍ���`�c���YY�.���K��!�=�V7?�ǥ'��C�GѶ�:z�]픘`���4ٕb��2Z���.`��7ҋ_gk�PW��FIQ�{�?./���@�A��]/ ��$�:��g�XK�2�O�@���0S���h��}n�&��G&�M|�2�A��F3r��KC?kp]~i{S6�/�^�~;I7��A���C���%��i��X���Lz���t0߿h�����.���r0��O�q�s�kkh�ٽ��'�S#~��rV%�|�0����U�� 56�w1Q�{g=����&��;��C���_�pj:�bf���|�e5�.5{�ۇ�����y>����X}�w��"����F�d㚗��.�_�"���J�u`�}ӄ�򹕔�����z�vP!�4�>�a��*flS^��=;)��U�6S%@�Ȍ�iE�3�X���=9�^�6��<>�c�
�GWY�,��#���"�EV_���;"��R���*v�k9��M\L �t�0a �s���`�f�3kk�i��*�z��??��&*�h)���^t��k�Ax��,+��nE�K�ElCJ*���C����N�Eg?���-�و�,Rf�6�^쭿x� 9�v����!K�X�����~��o���V�?rp���M�����V�\��<�rCn5��Mճ�	�d�4S��Ĩ@��k�o�[��Q�ݲBJ�g�f�JC�m8@x]B�x
�[�3���6ֿ7��A7�j,�{���4wU1�cd�wA?*c��d����x���%UM�3i9~��ƹ/�l�ߘ4R��>�D��@�MU�ts�HҢ�et	s��^O��f�G�|��c�-��ީ��g3��χ=�d;p��hz�QL�Z��g���Ig���ɼ�UXK�s��:H���,p�A0P{X�6�_ӖS��z�G�*���3�9��q����?�]R���r$q�0ְ�X�])�>��9������J��˥/��6�s������"o�[�� \7����5�BD���=ƪ((�[d����b� �-M���Vy\h���1K�#�"���i W�~6��3�Z��׿��Z��x�1|�����ݿ���9�������SȲ�6�����1A��B�k0KԦ��[D"�fw��J�u��<�<��1�S��,���^�W.y��v����]nf�r�5.�j65�ɾ�&f�`�݆ x��`��A6q9��g�: ��Qg��26��%����_/.�Y��ѧ�aP��Ki�#�S/|n��Hn�KY��3��ا{�XcY�v@���F��S�K6ۉ�G���y@b~a;X�N�ݬc����}���4�����z�h?�%��;7�-+�s[/��	53�m�O����2��d"u粎g�����jn{'���uPaQ����z���!6��9VA�m�) �ux�*�v�`���UƳ���� �ꄞ�Μt+;'�q�ԏ�x_?���zK���-�0��3{��s�3>���kKi`j(��F�q��p�"����,�]��Y*�~��N:���^�p���$j�+���w�������������(C��d����4ZǱ���wҶ|�1��� �vŶJ��r�Q���<����K����=��:aL�Ho5t4g��kߞ�E~<��N-�t��:� �1"!���{'�2'��@k-sr)��_��/���
䀐C8�8aD��"��t���Íb��=�� �7#��WV��7��lI������[^H�2��l����Pz�=���݆���&9:�&r�>�����mi*�g��I��yÛ:�%.t#K
l��}�0"wdvg�8A�ae��t���*)�	rb�����<!M�JH�o�J9�h��FgcϮ��:���EL���U�U�ji`s0s��e���Bܪ
��dV;���=�M6]pd2M��U�&�a�T��ğ��0v����|ԥ�i���#YαǯkJ�?۫ f�?�^��J��k7�3M�Y��w�@�Ds�G@��n-ڗ�52�[�2�c�xp{!)W��F�85��,B���f�� ��5L��X�}�z6*O`�d|�g� ��	w��x	�� �h�����'�I|�A1܅sx���8JG�x"�HL�@&����&�{b�؃Iv�Kw� 9_�nGZ����H6wG��;Xz
�L�ea�ST�y�֩�n� pK�l�ǆs1G�s�`�}�٫K����_����
7�ϫ��s��!�*�g�cG���~�����i3�e���q��HrEM3��6�Fg��Ż] �-���k���l/a�Z;���9L��WK�!�$��/|��P5.��\��/��j������?2�A�	�F�œLpi[rG�ps�zk���T�l&�l��=����/���MgO�-݆ m�\�a�B(�5�t�'nq73�9�����ax�h������y�9���u$݊ �O������۵#��ZSɛ�7G��47w�\aj�^��:�@�9�l6�7��nE��vOc_�r�a����Y�R�|��9�������B�_ 0�c�E��+�=��a}"�}]�N�7�=ĈdC}h�(���<�q��|�{��s���F�vT�?�N��,�7�g#��Q�A@���K���>�"����RV�Ɂ_�]v��cG�R0����#���/�J����=h �����3#���>GD/A�ck�e��m�^�΍Y�:CLЇ�`�J?�r�(��������2Ɂg������zg�����Ϸ������}��i�4}�m�t=��|��1WÓ���j��Qt=y�������o���(��%����RE� 5���M�\��/��Gj�������MŕM��oy�r[�h�ǌ��Y"Q��^X/�q�A���̭���:��P���#�NT1���@�*������8ŏt�[�݂ �I s{D�mf�&F����7�8�'�1�w43��vӣ��ТM�B��T\̞�(VOW��S���Í�3i����ޣ��sn7y��Z��9�#�O&�������b7���PA48}
��A���[@p�F���Ә0��:,��+p�r �έI~)d�u�.����\�T�P�������ۄ�.��N�q��ؖbz�]Yu�|]c�M�[]�BU�  ��J���=�i	-XcF��a1���H�]�-�8�'??��h}����p��,���AG���D�|���r,�[�R���:H� -���U���*%�*���v�Ev��Z`d#;��e�Q��"�&��9���ZI�!�pi�a�Z\@3�,��j
d�B>��a�4��|zB������d�E
\����w8`��a$�ɶ���\�".���b��3h�CqH�p�̮���t6�������Z:yTd�@�O,_,56�Frt�T��(7w	!A3�[���'
ܵ����[�bHk���9���^�fH�H;H���!h�Y�:-:h�Y���O1�&�����-��]#6p���N��T����K��Z���v��ң�mv�5��E�$�������=�qx���7��-��:� �#�_ĭ�t��{_�:{d��"\�I�����?a�C�S���{���<�ݬ]Y�"p MO���n���,K��Z���ܩi�w�+�[#���U:�A0�v��W��b�׮m"v|6=[%���ˎ�nG���G�!�D�NS���cU%�����R�j�.]
 �\�V��m9��%��b����.u���}�1|�mT�Ɠ�dZA�Z����(�I�t펻�T>[܄C���	��(�5L��9�@K(�b�?��cp�pv�#��s1G�T�g�y�9��Z��G	o�&v�3-s8��d8�~�ڡ���.�yc���v���% �kr����J�ꁋ�K��4Hd���rvՒ?�k4$���`�ǅ��3_l!����W_��n |(�!�Dk����Ȝ��ְ=�-�bvk^Y�(��v�g71:OTRQ*FQ,>2@�o1#%D"��֟�Ӈ玎����f���W��0�*z�	���L���1�M�%^� ��q��{��di�Gn
��e�+��aDF������#���Gz�7�ѿ��+�~)�B��?������������^t�|t{22�Qm�"K����k<�͟r��;G�4a�ě�s�W�z�Y���ޘ8\b"��*�W�l����O6KG�f��>�́���h���&�Gݥs1!2��8��M�;��X� �Qu�pYă5��5�X-��7����� �����okKDRjX�!�@:#��5�_�sA���]��ޜ_#�\ 	�}#��>˪s9����wfD�󧼵�����Ig�6�i�|���j���Gy���5Z�����\$9����ӻ��Y�%J���y�OF�z���+�\T0s4�����Q��Kˌ.v�A.�"]$�(GT�qԈ����vث�Cc%�|��kh3� CJ �����;�9��)F�Ҕ�r2��2<O��zD,-�DP��tb�P������T�u�Q^�?�/P��5 :���
��Yl�z�,�A�g�JZ��\^:�'gdl� ְ�p����H�3:�!������N�ggm����꩑?�D��w�b�ӡ��&}�������jN:Է�hT��t魂�ʨ�/D�3�#F��G�mF�>���I��a�A<v�w��DV� �?'d�.V��8rG��ff��<�f�x���#2�e�������R�:,Y�6
<%U��̗ۤN�ŎN��>G�9�3���>�(j݈@ـ @t:�!�,�eZXgWI�Fw}��SĪ���qՃF9
� �,5}�1/~�%����]"�H��b�&���R���!���YZ ����@��8A0,���4c�O�A�	���]u�,�N�Ztw3Ă<��co��XO7�j��1�?1�~rxR��o�=�APi�ӡ���eˌ��3�����	�ݎ�/�%s'ہw�x�ck�7V~��`�{��	��.؟���<��ی��/.�,T��0Rt}���;��Ϥ7ײAw�M��>}�[xt8s�ɟ��p�$5��#��q�{�ä����Dm�K(�v��q#D�!���x�nJ�]��R�H��;8��31�g	��W"�3��3�A�+��Ii�]T��=L����צ��5/�)�������x�G<���m�j��C<n:u���/��u,KF3�YN6��Z�ˎQq���nZn����㊤f���|Y�Z)A#�C�:��<{ڔ�:mr7F���e�»7G�*��eX���ס���O�T�4y~��/�z���nA  #9�f�9Z��p/�����Z�c����zҹG$˲b�f���jA���=�虫�H�����7��Z�u��x~�,�AB�ĥ�T�.;�ɲ3�*^H���g�N�h�Һ1�Б9�ֳ{�2��X����gFz���bg�����ea�'�G˪)�9����?�Z!���_�v������Kw�~w	mɯ�?�B����j��h���2*�Icw�ۓ�bWQ���K��Og�����Ӥ�zK �ʐ�B�2�J��Y��C{\t\:E���B�7�֋6�4֦` P����>����c�Of��Г%^��7�?,�.9��D�[��Y'�-z�\+�ḧ8!��u����㛣�Mh�A�\V\O��;kh����g�/"�_z��d@A6�C3���7��S֩��K�-DӘXO|���d�XÁF6��˃��t�t�`�4�ɯ ���j�ꆦ	�眱I��B����$^9�$Z�����¥#�z���K6�CY��@R5����۔��0u⅑��zO��K��-����S1j#ȸB�f�H;ђMe�2��&� U��#��� #���`~�Ȓ�R��1��*&�15s/��|���5 �ͥX��=N�8�}f�p����13���{P
Kj:�ćfl�q^ϓ8d�\ēޒWC��.��Nz07�d�d�~��tΣ����U�Z��o|mDШ� �p`��{��R �B��}��kN66���xXB���v�K�u�:7\~C�e�z8H�c���fA �.�Q#0�����
�Ce�
��nj�v����,5.H��@�����*��o���˾$H2N�����\��{>�HӮD��%@�u�,#��
����K��|B�6�A����^@�aƂ�ˎK�\����.C �>C��}�Bd5.6�9ad�H��wL?󿗳���[�#G�]��\T@ߑBC�y���A������7��J+��J�=_��/������ŵXn������+�Wb�ܻ��Ҟ��-��;�Y/+�n|e�t!�PR"fba��Q�~���W�
��^0s���ra;��
���I�I#4,��J&2慺������ב�i/��[\\^����m�A�XvP	���o�ѢZ��:���F�6R�^5��yn�gX��%���Uņ��C�FC���TcY\]��il25��Q��4cm���Z�nC�ݥ%d�iq�;���<�km��l�����G��Y��V��뼻���7<����������#�~������,·�?OiAu�7ۥ�{W�m�`w;2"����/\�?7���ƽ���4A@�~����2^��ueTT�����1;�^;Tv��5.�4܆�]�3Q�g	$�Lf$�+ ����"���%b�	��:����w��5�ה���;���%FЯkK�Q,w�&�`�t~�J��ﱛ�B�ltc�4���%�±�2���d�h9ֳ�B����l�����UG']Oqw,iv$ߝ����j}*�b�8����"�+",���\)�:�`f�qCb(�����/64+r/��u�A\�z�> �41:Pt.^o,�?"�*�Zh%s��5o�Z=�Xĺpm�D�Ϯ_���|1;ځ�H6���#��ݰG$
_M-��4�m̭���1z��H�X���c�X��W�t�v���~Ҷ��Hs#���@ri7��`��	�1��]p�Q�E*��q%��E�ŒDLb���ۄ� 6X�^����ϝ�[�ZR@j�%��pI�XD���A�g�:5�.;��$�n}c-�;6I~� �a�O��^[+����j��f�WE�	�o��#�zr���
{��PJǵ�;1���c�4UH�w��� ��*[�c�p��bI��p�"Z�-?���QgDa��s�.�!�a�唃����{Q-�_ՌdG����:��@+(���mo��,�/�pE6�t� 6hr���,Q���.�8i�kd�t���M6�7��^|�{Y޹<��4�l�J�����H����=�i���7��U�*T��[e��#�~�G���l'C��������d�41�cD
��E���s��h�d<����t���Z���w�eu�=W�^2P�k>��ۄ�M���BƂ,����5\�My��%�7Ѩ�3��(*��ђ�{@@Oð�X��.�Y�0�2���{`l���"�cl: �u��õz�����pD2M�z�hl�'��4b��pP��F�ع %M8�! �lA���?����D�×n���S��b�����Q�Þ��Ɉ��4�io�h=?Law�+/	U?ٽ�ןy�W�zl���#vr����R6sK��!r����_�ߢ������)
�����h:���UX��{��#,�_�sB;~�eGq=mʩ���SC�]���3Z�6���1����L���~���f����pP�5/�e��H�����MCٸc��x5��}F"�Ǌ[�2О�$���《7<N��]�B��S��������|��b;�:8`�jE�>�'��vz��ߗ�J�(!ih=��e{ե�቟3��tl������5�E�V�#1l�}���`�oIc�e\�����?��'��tl��6�'��NBX��5���mN���'��.�6`�7A��ړӤ����A4��Ϭ���Љ��혼�o�sĆ�Տ~5�-q?���`�1�D��^I���XҌ4�R�y�	N �wxgP-��"6�a��noX��k���_`X����X�`#4�~��%���8~'�n�q�@ҰL�4X�M{��F��u���Ng��T��rV7�Y1���]��v_[��Dz�`�g��],g�A� �����������,-���a1�4��}Xr���P�A�����1t�@J�fu�k��K��V4��w�f>>JX�Fk��КMh�gY�suW�.1�u��ѓ_�дˇ��C�9�i��C��WˎԾ?=>s;�p��pH2� �b/�Vn+��X���>(<��}c��s@J0��QC���E������{^�������щ�ey�A�#icn���ݯF�就+WO�Qߨr
�k��fm.�I/'PYc�On��i���F
�_E�,�ㆆP@l ���N���N���X,�=�	j�X�Z���:ix(s@8g��^��m��)�F�|l5��F�����-�AI�	������5Q"m���_F���Q�A4o��^��D�GG�1�BX�;��[(.����ep��).�n�N?��7���ڶt�PL���<:��$0$�6n4����=06��2�Y�z�)��Θ�|:��f��%�۶;�������'}����N�E�1���j�Pj����,�5���y;��M�/��e/�pF&���7QbH��'k�QSO����?�ߙJ3N���Q:�~�����M��^B���H�J1A���!�Q��>6};]<p���G�� ���쳕�Y�Z3�S8��r��C�bM8�6p����ӛ����ڶ�sd�t���|#�O����u~6M�M�8p�`f�l�Z����{�Y�tjF��ym���2��	����.�s����8��{�<������I�ȟ�x"G�ĶWF�/��yF�6p2X͝�ί|�aĦ�� �8�����9�W;8���DY��4T$�7�'�'���NcY�r��i6K�7���tA#�ii��;�Y�p�mf����&���%�N��*�������p�p��P�"���%��3��x��[���,|3(��&��%)a5_��
�+���30�X
�J���p�I�}��E�40��Rê?-�R8���������Kf��NP+�&�syzx��u�
g�{>��8���y)T���Ή'��`����\�'�⃝5������|αgéjh'�N_{����w��n8���ib8�0��w��J/8^�A������Q�ē�P�Em�?OrCi4��ZZYO���W6;�����|lLsߺ�8!(�D���uf8�3�>]_C�s�$Ґ�����3pb������������k�3-����Z�����3�F&�e8�f8�2��2<pBi �in��3��<g���v������x��3k4?�/�Y�sU8!��<�׿�'?p`ÎO����s�sK�=���;,�O8��bd�� pq1�`�F��b�3�n@�+oz�|t2ճ(2��'��lc����C`���n8�D�_��q���m�3�ez���1��ڐ������g��yP8!�p\<�/0\{�L�K�l.��cd|�F�3\��p2�p��Lp�fX>��<p���v[��ظ�a���C&8�<�P��6pv�Z]t9ù���PM�?M�sڒW��?B����X�|����o� �4n�m���� ײ��U5�;��u#s��N�?��Ͳ���� j(�2����,����j~y��%�8^��MSgp��v�wx/�����1�B�+i�/:_�{�	��=ӿ1�U	�h0�k�קѷY�Χ��2�����5��=��� �,6��(梭��e{�VO��ڨWD�H�L��W�v�#�n80ְ!�ŏ���x��s��pb���&�S0����3 �#��pl,��κ�'O#+��^�g�)�`8����`�8!+#��ŵz���cO�X3��f��/ȯe��ZR�N5Á$���XD��չ�u���'ng	*f�ls��<�A�pL�i?�7�
�653������W z���z��a[�Kn���hM�_���xw|1�fOˌȒ�@�3(�T�<�Z��C3W2�"XE��Ս�m�8��2���!�%"��>����nX�$p*�����@�i[�������`����f��o^�ڲf�M�	�GH\P=�w����#
���?�-���\B@zJ냂Bj'��Ia���� r����E|�H�,��b,Hq%��g��]~��|>��q)<#�����`�Yt�&8� n8�,-���d��L��p~b8�&82Q?���AL7�x��#�=����$31 ���_){`�p`���e�;���ہ�|:��q	<,�3��׆tgX\���h��3�y��,s�{���'���|/<�"��,��$>(A %��xW��7�����<���F�F�%���VoH���:�vXW�� g%{��Of7�'����.���h��{wguQ��q�)�7p��Ď�lbN��ء8k٣������	�*�F[p��d|�ء8�Kb���^t�n8�����lci��Ӹ��	����N�����( IS'�p{����6�ީ���b��v ��2��p$�鈋�7�8�tg9��|�t�u���Z���k���v����p�9���	���B5�?:�Hƻ����3�r�,��d��;�������_�/q1�x�<�%,�x �&�eq��3��sG�&8���DN':V��߯	�pz�� )��V0�s� gs��0��t�g)�s�-�t]�K"p 8}Lpv��8;��	�Z����ւ>.X��S<�XpT� 6�nD�����pY�{���y>��
�8�M��}]��a8V���8;X�|̰�
'��� Ə�[�lL�{���]�2���tr���|k\8��u!SW\b<ȁ!.��[�����/8༆��hOp@xS�Ϗa	)�=S>��ɲ����|���>NA�?�u�W�ko_@���E�p�'Dj
��@n���)��,��`��z    IEND�B`�PK   �C]YR9��b  �%  /   images/81a2be6c-b468-4131-a428-4eb848a41f07.png�z4�]ׯ�N���c���nB��im���-5���-��E��D=�.QBD�^�x�<��|w���~����u���/���o������Yk��`:��(((N��j]'?Q�MGC��*�ё�8]Ko�q;�eMA�p�1� Z("�n�p��q�Q_�j>88�M Ўw�rm#�A� �e%q�h'��m�3E�� !(��*@�G�L��&�>n��E�o�����n	 �7�E�q< �04hb�h DBJJJ�!�y��� HIJ�HH�K��@`)Ei�����$+ģ�k]�����t"q��������X���HHJIHI���ם���`�B�x��������'Q��
7ܟ��_�"�L��� �KJ�D!���<�)G!%Юh7�;�@Ƃ��✰D,�	�7����빸���&����M0�š%��	XO<��E���?į��W���?�����=�/F�}0=��S�ģ�D,��u�#|��p�� G�8".).	�r K��) �M ���:���Nx�Z�/|h-rSK�$! )S)iEYEi򧌢���PC,
���O������B�q�����B*:`�np�a���h	��#���+jb]�x�b2��oԆ��z�"����R�{�1��)���� ��
$��!��� 9BA,	�B��!��Ez����"���
G�e!(9I��)�e� �\��H�Q�(--��5<�\�e=��̈B���H$�����)�g%-�)ȁ�R2R��r�d���ᘆ,?N? �W��qT�z��HI�/	�������1~�Cv�pP��Մ\�Ȏ�������o��A�ZhaȖ~#���u��/C
�����w7�b���ULL���\1��RP��}����Ս�'���s����Nh����X�7��p${�?M���� ��ז!�r�
(0�N2 yiG���
2H� �����5w�/X���wwD�7:���V4XZNN���8H���p�<�"'����XZ��[�Xw/4�/Q������'� �t ԯ��rG�Q�q�(
� b��m���c����?�����k��+������?J���\�~��ߝ|�؍�m��Q�ˣ��������t�������"�
��'R�ǟgZ�;�ox򉵧#y���;AOK��'uɖ��t�^�uM���v��(����i��SU�[ذ[�\d�����>0�tɿ��Ŷ0p=ڪ xF�Q[� +?���?.���c� ��`�i���|�+vY*Aɻ{|�;Xi.��F��5��5��.���� ^����hUc#��I�)��m� <̑u��P]����p�*^@'��;����i����'q"���_e�㓨����鶢�x�5������ǮI�7ٞpI��i��:3q�Zpv�	�7S#���f`h�1�'�~-̬3�,_c���.w�/n0*R:����H��y�mSo�f�L�`Ee�����p�9k��ׯ�B�Ņ��k|�5���Sꔳ�ț���dzf՚�%���'j�����!��2��ݨӗ`QSo"k��HF�1�o�Y"�f��Qn{�=8�Lx���fE��ɦҐ�|��B��սwF�-`����W�޷��;�v��(�&��V�vO)zWk��kqw�Pݵ�C`���;�Y�m��� #���/Y\��5���9�+]�-v5�
��HQ�s���vT��>���x�~��߀YP�u��2����F�����4�\��-u�+\����L�bBB�^L�ItY4��Ǐ��.D	�ų�� 0EJOP�������QuQ	���a񒧧�_�kv�=^����ٯ���LV��2o�8=����e�*z�w]4���Sy��V�k}��xk���"8=?35�F����²��p����L[a�'X}��2�̮��4%o�n��y���u��R)���aw�K���g��K��Ħ�R�y��	�I
�˒�ݹ�8!++{��s�[���$9������'@=-�2�b%��'���a��R����ƳC���k�2�'�;�����p1ۣP��� ��.�[ν��~c|���}dp'[;����@�wG�O�{D*��|�������c�e�㮡�u�!ȝ0|F�!k�hd?gK�&T���L@X�e��Jv���
D'����Ť�$��2���C�	�އ��j�����c�S���d��P)ߜl^�Sڔ=_G6N��;�y������yRy�uuʧ�H�7�Q�}�<i�ÚĐ�֟�P��sx���A���L��6�)���s6O55=P0g|k@xB�����fm�5�ID�
���h�EҰ�4_���h'\nU,ʿ<��#wū�1��:S��Y$=:-�\����/��(���gLF��g��e}Nb����Z^����"n���K���T����ȼӔp'V��;F��^a�M��� ʣAT�+���U�t�]n")X*�D7��Uk�9����B�0��#�� �|{&�����ݫ&	šK�ؠ®�WW�S�[8�"+x�K�����@]�������cnm�vRE�p��P*�l�7��J�_P���y�S��l9ADy�(wC�v �Kr妶�#�Y�{��0�	��Oy'2e[�C��D����g
�x�E�q��,�;���)Ŧ[v���V��jYm a��\n_����{�+�8�l���{���R'��Je�,�t�I���_j�űH�O|ܠ��L���4���Sc�<��{5<KF���~�#*H�]�Pl�/�ͪ����C�.�0�a��M��^{`�CWyn��bZ3$W�^ѥ�d�T�xo@?���������o��C��2�����T�x�㠕�1������:�����G���%u����V�4]�o�3�	_;�kU�Z�"}˩W�	�C��.�&��^ۀf��97����HL���(��@ݓ����E"?o�+�������9��7S1��������f��k�l;�U�»��w�L��<�|w3��%&�5r�(�� ��57xO�^���%�/�b
M�%���;��҉��;�=~��l�Kp�k,�*� �}Z�sn%w6W��{�f�6�{���Eabw�|���⺒zu�'L:�ʚ�mS�xe����@�CX��'����M���m��p��~b���s�V��������@HkYZ�AǏ��ف:r����(IAf����
�����r{������E�!��U�s��2��O�{�:�X||U�xA�j��ܗYV���7+�.7:��A�a�ь�ͻ�^G�C�@Qя��a߸)�l>�V`c���6Xү��r:��7�Z�r�sh�}
׉Oc�]6e�}S%M	��7��?Έ;�isE�2���ɻ��:��'�wR�i&W|TD}�JDr}9u��m�fr�ٗ�А��T��t�Et_�@u�x�TIL���C���ы,a)3Q�I�L��=�7?Nu|0�μb�=��h�|�3���%W��O������9��"�/�wr}
سۀ�q��Z���?�`������bH+�K,+"��\}�>���[t�]hv����67�o8.�˭��G-�q�*t���z?��t}(�+55���үy���x�>7��%?x/e��d�Q5�Pq��ߚM��h�O�@��h�jPM=�8E��$B���n���dIL�C�����9���m��DSQ7�h���]]���G���ym浩��!c�й�id}QJJ��j�v�^*<�0�r��unR_?<���s�t��K�q��|�b��񬪰��"w�U&���-�/�t��zb)C.m��n<|h��T��z&��qZ��%�I?��u����r_�P�R}v�~��O��[��{�5#�G;��~\�I��TB����hYe�;��߽;��޿5�i!�-�R6z�MU���'*)��}rZMb�;��1-ޓ"�l�ҥM{%*����y-1�DroG4���l���ss�����θ/m�)�wM]���a ^3(yv��V�ڸ�P%>�cǺv���I�5��kh�eDPfm*����>:��MT��Sip��h�nI�w�lvE����皊3c����_]J�i�ǳ�y��54#N�h�K�A_=I1'�i�������a�T�Bp��N+~�z���2?����>xp��
�����6��{��toS�o���SѬ�ԞUU=��P뵩k�!G{������}y��D͢VO_�r�(D2�f�>!J]�\4[��Xz��}�^'�n��є�����=��l�Zά���uƝ=|����]�->C�F����.
}�Bzxy�g��N2M�qD�ˑ�����,G4��y����:#�j"������P�y�����-�B8b����w�ei ��.Ǩה*��(�����a)K��|�Bt��0	I�_�k��QG�*����;m]lm�!��t�T��.�g�M�:Ӕ=�2dD��UB��'���(�.U/,0�������F2��ȇQ�� ����`�M�si��eR�$&�8�?$��|H������V���ϽF��*4�������by�-c��a4��9ؽ����o�b�z+�s
F��=����}��KØ�W���M	�Eu����},��Ͷ���Լ��)	�p���ɏ��IN��xZ��Ґ���p9�]��s��p�ff��T�����`nY�u��G��-��_�u�|�aE���ۖ��F˩�p�:͈�������u�i�UI\A��b�����MlX��}���a�Hc3 R@u�F]��m�-��3�jWm��{X���OP:�������.��#�T�Z�������q]t=a�Z�`P@zccc1s�g����oֹ��Ү�^�Y	"4���1oh�3ȇ�iJ9�ݑ�뭦��������xms�h��uP*k~��Y�j����w�I�&� iE����l�3g��z��v�}� !i���\=�TO��,��!���7���(��i�"U+�����&�^`]T�Ѳ�n��L��=
�|N�33�����������~�m��Dk��/{˷��kKJ.���O�n̥j��`�n���RR"�^�t�m	R���/O�0ˎA���z�,u6�yT�}����q8a�uɩ�q;�'s�v}��
��]V{��P�����[�7��^\s����΄��u�߾0`|�j[�ø�IV�c��ى ��ш	�~�s�4�E�_q|��ʖ�[z�43h��ڵ��h$e��Yd�H�|�@۩Ce� ^h�QBm5��ߪ�Z쥖�rz佀Ֆ5��F�*��(�:~����#�'窚��*&�sճtzS˽o.�2|��4e+�`]��d���t̸ĕ��(��qzN��L��N��I�,4%Q��Ml%���l�J��mh��"�Ð���
@���fC!��{`:���䑵﷜���{y���r:V����#۷�����
�NF��2����c��TJzј��5��a�˩oM�h��q�Vl�MJ�6</#:��m~�L�a��Sy[�:�R��9�b���}�����FoO���p:�>-*�G�ʎ.�!�O��sj.<y�b�}��yTi�Y��_��;/�sp��d�~�L.�����y^DR��ʥm/7'j6�g�����8�)��o�%X،$�A��������D5?��y���)��kq�Vj����T�W(t�V�Au�)!:��k�����B\Z��i�\
/�Pn�*̞����9�a}�'�
�8��.ʚ�izj$ކ6lُ2r[��C2B�	��+�T���.3����TTz��HL�M),�3��˻�E7����R��Q�b�^Z4�>����*���h�N,��\ߧ��&���h݀�QY�l�~V~g��w�Y�������^�d�gk�����+#�$m�<��bD�F;��U���J�_�"ag�cs��ѽf�Rk>�Py�'M��Y���jAb�mӈ<���6���F�jWEa�hA�V*���Q|>����ˊ� ВI�n��)�8�\�����(�1�Y�p��6{��;�UY���q��SLl�}#
/Ƣ'��5��AY-vͧm0B�w��<�/e�f���=�%.
��2��'�tX�����ҋ�
E�'u���.y�5Y9�GS���'LZ�����9K�ƕnQ��xc'xhN��Ii���ς��>9B������n[���q
���q��&��ʶ�B_���G-!'7�hXġc�.Î�d�	����n����-�U}��w3X�������1�N;��d΍]��`��~���rdĚ?�|Jʇܑ�F+��&J6�s�����P���9�~Z&n���R�~6�^����=�J�Q؈����!x���M��tx�A��@g��P2��2+��\^�<���?-�])�{>n&���i���(�d�j�I��i��j˩�d�`i~x^���SD��F��!l9����$�ֲM,��#�Zt��讌�w����~���7�b���ʩ_��q���;����~��g��Q~h���ر�1�e������B�a�r�S����p��آ[���׎�@$	�o�p���k�|�r�:#U̯`�W�{������e����ɕ��K�k�`��@�-���ƌ ������,4���k�3�����(;��G�X[��5IT[��!��q���A�gՂ��C&y ��n,���07=�h�Yn���xԚp��7��m�r^K��GT��ߓ���=��?�����ܿ�#�<�=���c/wݾ���'�{���z�܊7^����vE�|�Vjx~�.�G,T-��ҧ�s8�r|&h��0[sO�����`�Y�mNk�𫁊Y\g��&X��V���s�!�:=��ó��x��r��[��,�W�Aw:X�v�W �X@�m7;�����o4��E�f��H8x�TzZS�x�����9�� �@n#�/F�P���%����'� ��6���g�0��).���ٛy/*b�1���#�b%I�a��1�M@"�B���_��V���9!��X?�x�˗��p�9������k7F�i�Fb5y�W*9t�[�1��݇l��1^]B���W���wdA�y�08U}G�R���
hh�XJ�]�~m�jqqaܙ(o�39/��@ �l��)[�$%m+��(Z�UR6+�1lYh�?w�w�U�Y^�F���Q��B������-�-��Ѿʽ�o��-���.����߰�އIbH��`��uRTT�_����M��{�vk�1ӄ!�/�%��Л-=��瀂!�����ɝӪ��e�=<<G^z��S�\���E����AF\���oO@[�8�}n�7����3bn6������BX!I�l	���mH�P�#+?�!xoE�����X}��~M���֏F�>���(e��`xN�������H'5�U�S�����
�P)�X<�NMU��-�ˍ���3��0V���X�M�,W��#������5i��s�w掭 ,��s���6MJX�h�+B5��Bq�\_p>'��p�ɖ����xa�}�Ƿ͘�S[�K��Y_�L|��d���u�/��6�*+%$�B^���M}h� ���n�P�[��ϗ;I ����lɯ�J���ϋ�����y��O��qq+�f,p(O,��ނ��* WGS�B�6�;\P���|���%���{=�}�_q椲Y���ú�ʹ��5M�$���e�jYx��'��?O9e�,Z��fǤe�0kY޻'��]&���F��p��7T�MHi�`~�T�m/����d��i^KNe��D�9,���<�F�\'�H��V��R�zQE����f|���&~Ĳz{�]���`!oB>� nbҿ�ϑ������O��`�.��{�f�b��*���6�[�g��K��]f� 	�o��d{�粛�`~�k����fF�y�Y���j^�p}h�$vF��Q�<�[�׶�������c������z��? PK   �F]Yd��  �   /   images/83c9e9de-0e54-4db6-8a4b-a33510724988.png�weS�$��������uq��5���]<���,w�{޺�r�n�z�����L��Dk�)����@AA�+)��c����e����J�JCA�'��Y��W#�(ݠ�Pq��PY9D����r�V��"�����0;�;7����+�סU���ept�����?Av.~.>~��m�6�3����PH�x���ĕ�y��=�o��W�X�f^P<ޡ|��������M6ēb��HF'g��\$j���';H��g�&��Dg� ��}&出���«���_��z��e�k�	7E"#R4�өǒߥхx�[�����x�Q57���0\7)����/Pč��NK��|��	�I��;��*E�Φ�m��r.�c=���V�)�T��w�Rq��Гf��T�/�X���Q7|E43��<�I�|�)���	 Eʑ�G�Ž8���U�0�׊"!q8�/��ܗ��X�7��7�Ub:�zWY@_�˷���O�������ɹ0�a���Z�Z���VQ�9����VAE�P���!=G9<����j�P��I���IX�K�_ �My�����#��f���$���J�����H�o�uO��ٵ̈́0Z	�����ogs�;�6�d�
����"�2nl%n%�nm���h�]h	�K���.�T��	ų�̛�"��b#S�9UQX<���}�iFj��	��wa� Pp�9 �@�6���m5ߴ��є����$xM}Q������� t��R���Y�����S��I#s�h��x�$F�ԉb�����ѱ^�
o�
��Y�Է��|��ȏ죥������s���G���hY��*�5�`F��u6mCF����g�B"���0E���
gΞQ���N%�W��C����Oe#TS��J��ϕ})�ٿ�	�ŞUɛd���g߹���uk�����,�qp�
b%/*��˹і������<W��m�M6'+���`Ƌ���r�8���Y�� ��5��h��qa�GR�Y EM`=��M_�3�WV��XC�d;�%J�mڿ��Ϸ������	QV�1Jx��񮕝q���W=G��|�������9�y2�/RV�d�k��}� ^�o+��;C&�|@,4׳t��a�]���§����őA״vBt��@_m7"���J��^��ᾚ)�o�rj48o~�8�g���m�R�1WX��E�V�WEFb��r�b�kT҉� ���_�-/jF��C���ן��¿	i�J$ɒ0�!����������R�f(����;�l1⪖2u��.��$e�o;�(~��*+�n�9Up���9�J�״�����jQ�H�G{g�]��0f���-�DZ���T+N�l��:r�>YԊ�>��(z���0�2e���^g��R�3@�ot_~zai2Lp���&�D��y��>�n~��U�;�gIƸ���������p�}Gw��N-S��`,o���^
��{���iN�-�G��{ ��@#=�PX(�x�Y�[f���ClU�c�$��B	��l��eY����+��. R�n������a�Z��6�(�`|M��9x�V�qQa��0��S?/R*��\�1� ���CG)���G��<V7]��mo�N����������'EB�rS�H9Q����m��j�JSc�\�9FnD�b�d=��'��
�Ґ۞ʷ��q��ASG�Ơ��n,/�J��X�������`�D�;\��i��>�+�k���j�� Ǡ_����Dpb`W�~��LK|z9��K)���!!�9�s��(���0�$/�͵�g;�ۊ�p�@�� �orT/#� ��R����*R�E����Hc�J$���V�N�eև��:7�����>��a�������U+�1��P`OV�N�f�T,�@��:�=��7�!��"�Z:����̿�ᗶ�#-�P���͉�k5a ��9��r�ۈ��ft�!���0B��u��^2��0м��E�����Df�t�`Zw\����װ��jz����������Q�|�Xh���r� 3]����`ـ+��XEɇ��0B;�y���Xa�_��P�X�t9�W����'����	���"��-�:a,PV`m��3��8وf�#w��Ţ�
P��M��l{��A�{[崵x5YE yR�����@�>����q���H�'ԁ�U�� [�M0�DT��8ުW&�� ͳBd��aK��4�lʍc�1:S�ϋ�Y�������x0�W_LHHp�d���w�4�E���&�/+[QN����$�t��O�ŊE��L7��Y������՛+2�qW�JHȪ]WI�v�SBvw�'ů��D�&96a�H��+_к����/��]̦�\&~�J��y$���"����,����T�L�F6��׬���_q1����}P[�M,�~�'�(P�	���^�B�Bdv��V݋Ul���5�.Tt�5:L�~����d�<`[rW5��A�\��[�l%�m2�7='S;�ܘ�׀v�1B0��{�����O��(�wTN���Y����[��s"�@�tO�M��r�F]��9(����gj�1�k��	�g�
/f���G�@M��*��P�G3'�oK-��	���(�W,yUN��lF&��V�\T+jf�n2���$�G�b�D�.u~�N f,�6=� �E>c�h�J� �^�AD�Pß��%�0��Vє���X�Ђ���s.��j| ˈ�O{���q��01�5�UqI)��g0s�^;b)T��jku&��'=y��x�>�:�h��|a� ڎ����_�~��g[�L��&j��it`��%3�E�s!�I��R�=̣A����O��($t+�àɀ�)-uWX�dUU�[BdHD�"�e��,۞�e�������ft�o��x^h�v��t��[�"/k�ր�V�x�T*xJdy���EeϱÏ�ePi�Z�ZPg�3��^qK��״��4�f��4��Ua�ʻ��u���1�}1Z��f~g�ȴsg����Ӌ�~n�e���P]gSzW�ܡE�^�i�k*i�=�Hk�Â�AH�IHG8v�t�$"��"Z^����J��ȥ%S%v��_Ah�A�A穸A�d�DE����X��1�
���< ���~
3�'�R&��Y��/����C?�Z���2�Ws�|�nݪ!KR�N�����>�o���e��@,ŴQ�o��e,m φ���ߩ�Ȯ�D���˔�������K��o]ӵ�᤿��$����p�����؜���55�)����q�����ĚD�*��'�s�O>�4��B�&�~w��!Mp�a���:d4��S�q:�r������h$M��_�9��#,ik7���JZ�G�B󑷂�hVf��O�)�&���ګ��|<]���I$�8��lM�N֙���Y���@��_��B���epWq�D�Ē�XX31��fE�;*�&lO]��7,�%lh/
��ڭf����X��Ѝ�s������ޢ�4�P�)h,@���
:Hׯ!Ll�?���
,�'C^vI6��i�*i�M�GU�R�݉�1��G�c�~�Q�K�m�hm��V�	2�T�~O+��	mC�'`h B7��b��`��[���\���)e�24�+:�gH#�Z����.u���b,`�b�9{3�FH/@��N�gj��[��3�v��n6 Xߛ�k
Ƕ~?���op���y�@���Xh���%�����ZNY�iE��*c4���+�ZCڈki��y�nJ{sc��<hVp�l�B���� !.�m�Ӱ1Ei������K�Gk@�q�/FY�4�T��Tܙ��Z�1L�W���nc�U^q� Z�pӈÁ���X�{����:���H��q��M�ԭ����Zʠ7��&G{K�qU���.��*\�T��/x���؉� �*:mv8ȡ�m�Q���[Uy�^�n�<�Oъ�����7�_Mi�Gv��@VJ;X5�}w�c4+��h��#�%��^�<,��e,��i�F��8&���e�v?D��������br�=I�n��9s�*�/e�����.et�Ϋ��(���O#��2N9�&���ɫ8M�����Uψ���ƨ�E������x��n���6�e����Z�K�f���p�Y�|�Qp�DC���� �X�E����+�N �����t���Ka�T�xޚ�|���O�(ͥ��mY7'�XQ�m�&Y�A�������d���I� �n:e-���<2�q
�δ�傶o
ߌ��b�{���U�I0���ӟA[�VW� ��f!��l$(4�@��r�Sن#㡴b��]&AP�x��pb�
W���A�9��(V3b˲���apUIq�:֥E�]�ՈW-/|S��C
X�ԏ��oa���M�^a�ϠZǶ�T�k$���c��e�T!��e�����%W�����:v���1��G��iQ
SY�cb��hI��}FX��4��:��%-�{I����%?ϙV�77�U(.�W��g�¾Ά��S|���hs�u05F�阑����
5>�_�4�:�c�dF'<w��a���ߺzv�;�ZyV>E�Kb��9污T��Ҥߑ��t� $��n:��F�o�nd�}��ι��rڠ]W�ϵ���ROU�^��76e��?s ,����!���"�6���W� _�TT�����fj�o B��?`d���C�����\ҿ��L�9m�Y+z���ѳ�F�GV�oq㿓+J$�-�{I��5��-4��+փ�-�`j�\mP =�O#l���B����ڶ����i�w ���_��i�_%um�!�I��oq����*�Z^��m+����>�}ע>-5�e8�<�ITa6��d�<�I�-��5?�a��5�1f�g�zZvÕ�5�AцX*y��i�-:c]ys�a6�VY��i��{k�&3J�C�+zcW\`=�ך�n��fa�C�Ql��Q�^��RLE�L��83I)��&YrL��O�0i�q���kL��p'��y�������O����V���[��e�j�����[Ǧ�V�FB��1뇙_0�I��?f�y'�O���&n+ 8	R~���ULH$���)�P���e�T"r��F�P+��4 W���}�eǻR�F.NK��@-�rᨴs[�1�w�Eg���|�ܐJ(-c�\N�M,iX�Om��VAeU�H���Yy�hv>����L-�X;�v��x��H����X����bZ��4)k��O	`�IJl��YܶD��y�/�|W��wp()���3�ݏ�{Q{`��Ș(I��+,���Wg�����|���$F(�3.4G����nKiM��Zڂ���ŮN�b	B�[�6��r�l�$�+z�6�!_���Ӫ�j�)[ݸiY ��詛"1J�}�]�m9�d`h k`*6{���Um3�J�����*�X<W����pȇ�	��N�!>nQ�˽�3<���@�2����E˦�`��S36�� I�O��'���:���U�B�����G��|f��a64�k��`��Μu��V�� ֆ��L���E��1�?@9�-Kl��d�s�n�r���ap0\!����X̀≨Q��t2Y]�͜�_s���cDO� �x�t�Bc	K�!���� ���53M5h�/X*iZ_�㛕2���rP^t�C&�|�uE�z�[^�Q�@�AL�q���G�o�fn)�T�P���'O~�H]�8��i��5n.�!�9%��,R��

�!�I,ik���Qc��!�����<���#��� j"���h�l��/i��q$�:���������K#����v!NM���.�z��?�g�n4G�TV���y�p�<q�b�/3"ߒO�m�$p˾��+�������t9{|�
j��;��_�$N?x�a�
��y'����Y��^c�w�����G/�ER��ة���$�,]�dP���$��zg��\[�����4��۱���GQM�|�����C��/b�Ϛ�.�%i�J99;�5H��	�h����U-���(��.���&W�!��w0���T���'�_4��pDw!5�����L$�ms/�vϔ�"���v q�������}�a�1q��Y��i��/�c��IOa*VjR�E�"wҹ�)Ȩ��J�Za�t4��N�Z%\�45��>�|���q���[��w6���t�N�L\.�c&)�S myyjt�2T��FV������M��#>N�x��fJO�G�k�]U�C���:��k9�eK8#&\:�	J���O7�5�4�̵-�H��N������������㠻�l�'O)[��q��_3���}s3��+��¯��?�a�ڱZӣ��)��}� � ��:�~e�QK�jK�9�E5�3�`RA�3n_}��}�xX2��ԶA��R�J��<t�D�|W�g�'�R����}�LP�_�� �3���AlP�*�U�oh-�2�qS����p�E��&��s^��D�%�Yfh�Hˊ��m	<���|��3g������$�#��5��?�v�R��f�'#R;��ĈyY�#և�P�wÃ]�q�[}AF*/�t�;��F8��I�M-Kh��
~�T ��`o�}���ơ���8�7*I9ɰ�T���l"����Xs�o��?�����~��Y��Z�*�+�-P>�l^��^���O� :���I�홶�ZbM�=���-o�F0��{��u��4qS����������g/tX����۞����_[*/�A�z?�"%n>$�RW��<$TМZ��)>g�I��砃h���$�T��!�vIm����\�|����/jJ���r�~�
�Ke�CA^��-��������\f����#-�̿;��V4ih���X��W�����B;�"z$�1THZ�"�½Ρ�^V�W��P�.z�0&<����lP%����T�V� I� 1rدs���2Ѻ��رkZ��+���̾�q��o�`5cF�/5��g�y	�k3�}Tt?�͈,n+"�h�91�#BF%HgF}��x�0ug��%Uy���f�����y?v^꛹�.L0T��q�%�(���w4jn�m}��).��sm�l�ۏ����F��3f����m^�){m
_�BW���uz�f�Dm�m��c�.c���O��E����f���qb1��}!ߥh���]�)��jS�3��Zж��3K�u~7�f�c�ɇ3}۔�_*�PI,O!��+&d�՜��������&��z�8���Ţ@��	�3�IF�Q}�o�z{{?��L�)�v�J� ���j"��K��f��mm�Ǡ�c�;���?%>�8M�n���FU(�Fn!:��2c\g�p8�����;�r&���Je��� �V�U6��q�}�_)!,������e��}g��|]��K0���y	|������@�n.�����!�ż�;��pK� �>V��<��E�_�ĵ�ݛ��P="*3�����mH�oB���Jn���Q����ýۀ���A�k�ێ���g�h�¶��tn�2�qot�������^�����@�Sy�h��ʎkb	yDm8�٫B�Ǭ���cZ?0,]�cV6�ސ���ٍ�מ� N��/��j����_��51�����;m���ֽ�A�Y���|	��0:]�7���,���	�K���y����
��e�"+��[�����l^x�?�������\fe����P�ۄ9=����?�}���z��2$ܳګ�K���[�b�-�yA�ۙ��=n�4͒��v/�=�����a���t3?�}@
�|�e�y����H�����vi*����+����ݧk��؋�>G`nN���Y�f�}�~�p�w�K��ܳQy�7��ӹ�J�@$;����c/�K�eʀ-�������O���c/��OR��VK�ี�'K�ьxd����~4`�/��+��P�S��1�_PK   �F]YN�v4	� m� /   images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.png�{eT]�����ˠ��Kp	 �Cpw$�%H ��'��Kpwܝ�y��_{���9s���vUݺ%OU߉��*��F�  0d4  j  � ��B:��Bt�R��`�H�oT=w �P����S�^�����t���6s�X�Y�Z�[8;�譅�(ʼ��u�����.q6�n5&��h��H��tҠ��_���o_���ݰj�9�j`@LT_�Z��d���BX��%����T�^�O?�ڻ������;�^�t��#{{Thm�+��j���J;�?��G,d���)���'eH8����%cG��q,%5'��O�N-J��dj, 4��v8?Y#�0Ӎ��?�`.�V��z1�O�������{W�8�^����ap4/~b^���P��^���}��@��-:P��:{1��ΑW LQQ���Z?���U>�Z���N�1C�]ɅS7�HM�3���?�Y0��sZ�ۅ'� ���%,҄nl!���wD���`G�b+��O�~������)����,�J��z Rɻ$�-�TR�*Q8=g��?�Ѵ�Y iEH$#'Iz�oY����+�a8=��b0ҟ�B�T��}��;5ʻ�;$"�;W�P��$⛩�4�_g�,�� (7?�Ɣx0@b��awr��`��1hdb�Ծr����Cq�Ӿή*�Ä�݋�q����LR��\�v�Bo�`�z�̐��I,���F�4�!�����!�
@�p3O�ij���0.����ZeE"�X�%<|)�ؤ!�`3�2����a�ƈH?��¸�$�� ؈�H�QGjC�T�ژ�B�`̄y�#����vm&��"��[B��IL����g"����RhY-��C	�
�I�H�VAt2�w
�Z5����얜����e���!V�?���>4���>*$��H՚�n�	�RBx3N�K�#�u��_�u�a$����8�d D��1�J3 7I�*E�ưdB�������ʠ�DJ�~7�S���yj�d,�8#V��K����������,�cʪ�c��C�������b��Z�8]| d���f���g���sj�=�� ��x��!�&1�r�Ӕ�`�co����#��&�Q2G	��~��^klQ�0>�s�5d g�B=�d�H?�JsVP���/�ama��&��?X5]�(b�Y���ӣ@��w���'�.�7igi੅�)0��VK��E�i*W]�Tu;=�,����?��7q.N�;�.��ڴ�[P�B�6��[T����*.E��ہ-��'_sI4�Ҡ����:���=8R���	*�+��t�}�k���7b����{��>҉"�T>CG����WV�Z�����Qʈ��^�	�?��9�̫P/H�"��w�Z�S�;WT�x�6��:��I�R��E���� W�}�}�{�*К�ì{6\m��%k5'u�A�lK������l�	u��4�x�J�r��
e"
��ו�+)�3�+�֔�OhԠЏǻ��qF
.�^�TȦ<�dJj�_y�8=r�v��g�E���0�ۆSkJY���{��u_�#��H
߾��92��8���� R�b~�4u1p�iF����".pP��j���{�<���ٿ��Pu��,���t�ڰ)կ����ݵ̷��xv�լ)���;f��h�N�y��?���=E,��&&���;�"j2y�0R�H���)d�����m ؉����3�.� �U���ցm�l'�2y�1����&T�70vႝU_�X*�X��ˁܟ룽�����<׋y(a�Bᇇ��|�է�/�Vē�'�)�o��@i�_Gx�����I�UeO�Tl��	j��#��Q�TӃkw���G�C�#�X�ƛ9����2 j����J�xQ�eC� H�X�f����t��tPԯw�A�n�r�7}���R��uNOǈŜ.�{����U��	��z��잤�a;��ب	��2;�<�U���[�0�6CZ�zP ��$�;�k���1�����-��&}��ܢ�}2Bsh�쫠R㥭=�?��65$꧲
�Ɏ"|��b��{����|���M��^�$�0 q�$"��Yo�Mp�+�ڊ2�#⫩�+�>�����J��t+��)�W<!��K<^�>�ې���YO=����Q�%�rpb�Q\G�vË}il�
;͕`N����Ml���`Q�昷�;��O�S̯��O��R�>�}�Jwɑ��mq^���Z��o
~p�EI�DŢ7��M�������SI��C�2�YWT�N�I���#��
O�1 H4��\ԶP��@�^bG�A6~/h�N�K��'����"��Uo3�0��i�ZI9V~�9�(�<�Yk!fӁ�4B��e���%�jכ'>�4��?Hĉؓ��8�tˣw|�AbH*:�I��-FѴ�����M��.�����`�(S>��H���ϳ�� 3�m�j�=�r��.��fm9�B���!�+�nc�x��#�*����k�S�B�������ug�.U��?_�}$J���wB�`\��PL%���17���/���[�YS>n� 0^C2 hs��Vw���/l|���!��}#Vs�s�㐻W25��G���c��޷Y���LU��P�&�:����-|ԩX�z�Z��WM;W���*l��@;���Mc���x-s�������k�*��}��Y`}��� Mx3B�CU��_�:������N�%��WO^��b�*�z�oə�h�B�cNE��<���½׷N_�}�������ڑ�)^���L27oL��Bj�q��Ǒ�9��=(�}���s���=��D��	.<G����ׅ�!�8��t�v;ń2��Dc{C�-Q�g&#SN���Ō��_ -M
�㘑8]U����N�˳6���/E�`�G��f�eG�q���0C���g��2��JY�!>r�D�]
���~Ӷ�$x�H��C$c�pG%�]��� ��,��q���=5�f)a���1h*k^��G� >�s�bQ�E^��J����1�uYL�:�
���'��s�!�9q?j6\(�x}��c��"_�[C?i<=���)�v�e�Uhy�Q~�g��
]������F+9F�8�FƐ,�D��觬�B�.�1	�?O�y(�D��y�Y��"�P\��<�[s����c�U��ߙ�*Z?�H3R�C*Q�����-ȁ���*7�HN���^gA�또�s�����`U�D�mɩ�V�-����i
z�8G0�U�d��;�H���X�95��YE�*�y�Ħd�{|ej2}�� ��Nd��tw�"t�h7���"(�2�c�G��ɩMb�jj�t#a�G�����A&��!�Ԧ'�b�l(��E��4&2;��l�(>T靳�.N �+�F�����U�;��}�mv^�2�vd�Ϋ�%���N~���d��\��U���=�����3��]b^~?++�����3�1���8���
�i����d�H�K��Ѝgb���I �5���ҷ}+.�
&��!�25���Ք&Fa�7�0@�_����}�"Nl+�q���/��&qY���G�5�?(*�5fvD)TP�J�S�Ȉ��PW<R#>Y���W�l����<+V �BE����֜w��]�/؛.��ׂ��{�K�ޤ� EO8[+��Ӽ� �)+��4ro���T��`!��'��%�յ�::� cc�ٙ�M8��g��J�t-���k�ja]�~9:�k�W����t�+��$�]C�3��i�޹��F��=E5�Smi�?�ib�3����<ȯw|�����^�|�^D�7��[�]]j޻K	$Á�P��&(�MT��"�6r%O	�|ԯǳ'
�7-���;_���κ�9ME)zJ��������Zc�T�������7P�Lʀ�DyP	\�Hw2ny��S���J@��E(r�e��Wɾ�����s�R����E��36:duǩ�bĖ�*��~���i���}��;`''œ�§��Ξ���{�5���ɶ�%�Aj��K6��rባ����t��A�x��9��{�i�tCk���D�ٍ���a]��Q��_L3��|�wϥ��[Pp@�G�2
>�ʁE��F>�N�\Tzq�Ҋ� ���#`Ax��<)h��N`\���A�6���ċA���.	��-UȈ������ἐG=-�|xȤ��9�����-�q��[�?�~�!�v�;���;M����O-���Ѐ��3�HM=q�/{!c�� `���|�ү�*OK��0M�t���"*����_,�U/�������/�NM@�n��_g5�7Pi-,3�$�J��z�#r���H�#�'&l�ΰ��D�8U����2i,����V��{#8pB%���eq}�쉻�� k:PJ�Q�C\��𙦟�
���F�=cI��lv&�^��Ɍ��~�Նc���D��m����fWr�P�*�Ƅ�&�L�+��'U��¼�sB_�:`�ɯ	���S>���/Y��cG�vK�O� 8���>|Q~	�頳����p�� �.�k:	z	g �Wq��5r��k���?(�k���R����z�����=�bR3u�%H'v��~����]��'cd��;��֭��G,(y�����U������AVc�m��}�Y!�\�uL��P�b�;�Lyr��Q�"�T:u?��$`���^	�]T���WF�����1�[�����1����l<}<$�i�@2u����`��5��ù�p�\RII #��Xe��i\N���j�X�k?k�R���]���^�pa�x63 ��IYd��HI��&��!vy�o��֩����,�]1���K�}�������8����J���7����j�������u���+��u�$v	���F�eo����J��G+�9\��c��_*q��>����w
��S]f���٪|���(h8Q�D^�:������E�'�e �?�7�e	Pn���I*6�|s�W%�B4s����E<���Ĩp�S�w)��:��@5��솢���YPH2U$�&hh��;���k!tv|c���+�s�h�u��"�]+g��w�TQp��̔�=��k6�>ǡ�k,!�+TEWY �%�b�[/̀�������2&ȍX�*uY� �z-��K�h)6/Q��1���)��Kbldӡ6˟�@ַ��� /�IHۺP�gO��,���|���M�LQ;��7��� ��ޙ�-�x���o����V(Y���ܿ���S�)���i�D��}lY��*6���괷�Ľr���x����.��2S�]k<����G!�u:������AD�8S:"�Y��||�'��O���,$�Z�6C	��X�HD��)}!Hvʉ�5�@C�p��p{b�ň�H|�
��B�}AlJS»k/���^���_��#��}G]�&�6uN+�o~^��0��mQ���G%��[�ö�����r�~��C5�������ͪu��ֻ��%Ց�:�����J��UD}�06��=�[���EjɊ7O�]�F���?��u�-ř��k�V����s���I�<x)q�`"��{J����a.|%=:Ol34��+T
��zK��sN��<���2��g3��6�a��м��� �T�/��s���:}o�G�AE�cQ����o��i��i�`#���\�&W�=�h�/.��قIR@�Z���<�m�ݢ }����15�\�h&fk]�A�ۧ~'�ڑ�CKn[����H�x���� �Q�|�����S$�%�M���bgu~/�@*�3�&�rQZ���HL}�G.,>�g���栊LB�'%e�ԡ`+���X{�(�N�9"��U�~�3�W��?v���"wYz�dρ��w�BJ�̅_�&�7����k��pxMnй�9te^+����@��e��ȕ�o��M��\x|�iW�A�S�'���N-�B#Iq�+K���oY��WeL��OMD��\�<?�nu�>�)��y,�Τa�>w�t
:q��� ���6����!)���c���Q+�u%��p�-��̀��{��#]�p�iI���Ϋ�cR��b�6��ѩ��!��b���O+�b^��|ޭ�PP����*�B|�b��H�{>��}�S��.�Ć�^>O���m��`G1a��HĬy[�LAL�:��V��u% me��P��Tw)%AF�(,��`M 1��^�>�D���-ə��,]���ȩP�Y7���u���C�6�9��4B���>IƐE�v�;'H��2�.��+����j^���;cZ]�Łb�c�;�"��UT��G9������ij.T5�����'����j��k�98bu��o�"���ۮ��RLb@����Qv���,�$pCJ};x7�	6SN%�=�jw����$Z�h�t+��S�̇B/u�B�R�9��2��W9�t�t�.�TJx����)�6^�Q�;Z�i�%��͗e�m��1D��ߧ���ı���y	����#��px[I �� y������)$��4��8��-q�5�=fHz�z@�� �z;����#�ȫ�����jNF��K�I��7�)S�K�V��#���?�?�[����R>����g��9# g�'�~��_jZ;�V@1h�I7�?X��֧��H�Sr کh���*��"�Gb��\T
B���Pq����gek_��x�9�q���H<�iV^�~�_)�B�E�ANW�A�ːKU(N��Z�ﳂ�L
,�[5���P�Sr��N�Twʇ�[sq��D�λ��Ռ�0�����y^���Þ���4���T��U�h���w����>�{�[�c��W!@j�476�B��m�  �t�w�:�G�@B�&��TVXk�ͥr/��F�jВ�*�꩝>o�^�=PiN�cP�U^$�H��M����y������'8��ى��\k�W)�rw�~��+�(��K(ݸ�[��Ҫ��rYĄ�ԡ�&p��E���?άٝ�55��`�4=���O�hÞ���ϛ����лe?�K����/���M��,h�qB�w��5�oT��e�mq���8���k�j�`����BVU�3��e��e���C4�N8��&��p��+�Nd�Y���1��F�]�b��Q8g`}��lAx=,�AHng;Y>����G�Ga�5a��9jh֞�"���ڌ�bl�Es����rЮ�v�i��ٓ6�f��k�Qk�O҈���J'=�)8��Ԗ�.&n��y��&P�E����mc��]Z���x �~sc4���K�+0�LA�iz��Y��`|<���S^K��48�% �%���k,R�7&s�vx����)X
X��8��0D
�B�§���͈,ݒ��\P�T���R��I�`�U���i[`H"@=����S����}�q�=7�胵Fө�_�bo0kF�2���}u�ΘɁ~�G�B��6+��o�́sA�	.H� �|����"�k���;CRu�'�\��7G���
��#����Z�g~[��J�gyq6h��;�æ>�T}c��#�b��ێ�t��jɜ勷R�}���w��o��%s�`#�_�*J�u�>��us�P<[��#��X݄�Ћ��?��ce�G>vX&|A�1��-�!R��6,Pء��a8U�yY���ܡ�0ֈ�B3Ay��F�F�.ۣ�!����U�`��� 0`�W�Z� R�%ġ���孥8R�r���ͣ���E�����e�[4���؄~۰����/��]��f6�Nh��a���B<S�ݺ��z���w)�ЦgOսQ�!�hkN�ܨ����1�.���h�5���U�w4I-��7w}�(���sz����L�=!���r�Jf�å"xTe+^U�)�c��VcY��\O! �G�G�ZpDYY	��G�>�إD럜]�/���4�Z�\����UQa�i��_�F�B�Ǿ���$~FzXgв:����?�hU�J��#�`��YSk[�Ys���!�o�ꇻ��Џ{@T.)IU �|���g�~/��ij�Z@�iK� ��҅M��X�"M ��$&�o�O�1�8�*�܎��9% 1Fi��5Ź����qҹѻ �I���'��u<لc�- . �K��1I~Ħ.�A��?{�0�e�/��������qv�� H�4���v���Q��YHO�����`!Pe��'��st��^�^����GQ�����L�9Ro.��~�^�T@Ot���qrDـ�[6F&��j_ܜc�����P=l3�.���a���A�]E+�dN��޼�w�*�y��`�t�I"Y�v�W��Hhv��%�Ĳ�������-"�/ߡ{�A�b�%>Lfd�C|^f��]F��V�OB�/�U��,�:{L��k˂���W:@�7:���PÖ9�}�h<��@�6,u���F;M���[鈈d��H���m��Yq3��Ж jȣ�����+����ێ+�p�&�_�M[�(o����@G�=-�d�U�����*�pu����h��XV֦�4E���)���8ڮ���[.I�kdP��J��<�~b���k %x��{���v݅��\�~�(�\���;+�j�ix�;_�8o&���FK��� .3کB<�W�-һ�t� 6o�p1�i��޷�g��>�Fw�<\�>z�Z+G���s�|�|�e��Q�z�����{F�=����0m�B05�<�$���k��t�8����m[�%uY
l�$����J���� �u]B$i4Ch�E�1��]�_эCf�lcs�6�#\��%Ej�b���cQ��he(,�=��	�����1O37Ḻ��Yy|��wмE����V䤑�t��N0�a�J3?�������q8蓻֫��v\;��mE��0�H��?��-X{��
�����b�]@OB�����~���d�QLu�>X�f�����P���J~F��B-6��[��#]߳�1�oRl+|Y�o$�O�4��?
��J��������9�B�$���ʯ��V���F�Cɬh�4Pf�ϵ� ��D8�<�܄E{�;�k�]��e��d�A%`�=No�#ɉ��/6@#_��O]���4���(���F��Z0�Q��[ZwIss�d�O �)Ӿw��}bn1"�{vxwU��ŷ� (A_�i�#�m�������ӣ�ϲ'b���v�Iv�^N�ޘci@rM,�#n&s���6&w{'8a��{�Z*�/tAH%-q�,�h����϶�x���󚹯ߍ����#��=J��}Ύg³%F�zo'rC����U�d|$��V^�N����_��ZJ=��=�KlZ1�]r��?vtXc��OqYh1�e�:n��8�I���\Hi�.�{�9���[�NS<���w��o�ꮎ��Vۼ[3����R�?��\!�[8-bw�D����C���_���;huǼq������ro�C;F5��Ng���V�.|�"�D(\�ߧ�u���� H��y��1r<��Rֆ�]�֞��k�T�s�X�YRgU_ʡje�QX-� �4-#��u0J��+ɮC/(>�G�6a-4h˳F��o猙sՐ��ǒ9u�X'+&]�!��K%��~��},�m��"*�����c�·f*1u�ۭ�oo��}���yT��0"%�T�~�]��
��VTdÞ�(!@��k���1{�<��,��rY�5�=�
�V���l�U��"��E:����H���z绡1�w�N4ܵ��"�f��?���=�7�{6��*��D����VZI<U���i�s�W�3�c�ck���*�6]>�7!E?b�3ސ�d�lV���&x'�Y"�fQo��;W��۝�[<�em�y�&��/ʸ��'q��%���I���6���;������r�d����I3���^K��i^&�ԇ�o(�D�{Q~@e��W�*�	���)���D|����o��uQ�D.
��"��\ԁ��큮��[�1IA
���v�� :���<F�$�I�h���S�(��Y�M��Մ<��F,��\�g��ݒo��T.����w߄�LZ^U��5��c�w�
�DN�E��������A;Đ���>�����s��t��c�]q�>p�!aV�U`a0�b�v,�m:v�ٻ����軱W�������n���|�Z^�^���_�t�/���E��`��N��׎��؞_r��j���v�2?bŠ�D�u�� ѐDV�*a���!m�i���L�H��!�a3��/���ߓ�k�;(`W+ k���K��ETѿyv�����P��`���}+暘7<Ѩye�cS����P��*�$E���Cμ������\��ߙX��K+�*�0ȅ0C�s�V���'����J)f������4�՝~& J�جcILZ����6ɲ��H�Z�qD��4[�,�����Q:�iN�z�A�n�=�3e��4����m���?b=8�P�w���=Zl�E��$�ܮ��=��y=.5�/���6��b�J��#?ʀjN��ϳ�?���ęт3����ƨ��c�Ҳ��dL���HĜ��l�9Gۙs+*�8��a8Z��\8}�)�o�&`�r�R�	?n2�dWR�{�|Ya�Gr)|�Y>u��^��+YK�b,-���i�gRj<�{����]8���#�~�=� -��V�T�����8=3̴�.;��U:�;;�n�ii7%���Cд6�xʶ���m]���%T�]�����������b��":O�JV~/�^����=qЂн��	�Ш��olii;%�o�VVb��O���}n����=�Hcy��24ifap��B<���y��m��5/���v�5E�Egݾ�~��Ǔ���Ӣf�����{�&�Iz��N!T���0�|�${�Ϧ�w�`tŹ�pB�����4n�5��W�
C.2��r �s��Ɇ`0�JW�:rajo��E"���ÃR��B���=G���'Ku�ʋP�!s쳚8�J�P��>����Z{4�?6�[�{8V�����P�FVRTt�������y���5�ʲ�^1&HĞ���E}�-I�;,��A�S�%�P��U��v������M����d�D����%�	��k_�:{��TAoz�;�j�2 �����NB�w�O��lx2�Gd��1���b�A���H���]<Rw�>��#%|�����&O��D��|!f�ц���&gٸ扄f~�_�K�j������6Zy���:����̝Ij3�M�ojz|��b��6�P
�5c���a�}:�ڣ&��=qdiS��Ew'?�߅�>|�g"ͺ��n�Đ����U�� �ꚴk	�y���.]�^ň�������k��5t���(�ѝ2��4G�]�8xBa��2�7����<_Z|���ҍ1�;��u�n���}k��rU?�\�r�����ҍ�8<�/���7�7Z�M�G�$_3E�����N� A������hu���u�Z�K��̥fb�F�Qe��lk7�Y�7�[+!��u8����,�Wi�
i�h���Y~B�ţZ�F���N��@�}�/�o�րN-��aG��)��.ua���mRwҿ_��ϊSURrV�^�G�o�AB��~.���,J��vtk�ɛ�Ƿ�ht�ݦ�����ꕃ�c��6�H�M���\L ~�C�b����_C'C}ɤ:�W��TۺW�8�����A=k���#\��d�O�+9P��}�����?�{��D  I�iO0-�n/aX��׶~]>u�keo�H��B} ��ͳ4�Z��l��)@�5��.���I�M����
^,�q(��Bc���?�);�cOkQ1��x7��8W	5��/�&҅l�9|��:��?j�Ǧ[TpW"x��/}v��w)�����9��������썿Ͱ��qp�h���)!�="/ap�.5��GL��(�V�ty�O�{&�)J!ֆ��7=Y�V̧���MH���:��|A��0�+�vq�pM{O����Q�w��t	�]kr,��6�C��3c�ɑ˷�l=9e�㟔�}u�A��R�ѦZ�ˈ�[�_�#Օ��u��xw(�\,=::��m�h���)!qk<"�ی�/��.;�O�2ȏ���Y_�~U��~�}�ҹ j>�K��&�v���X�1�����w������g��J���������67�-�k��$)!y!c�?��7����9
�����]�����C�	j�����{
R/��]}�
�Y���K�^Y�y�5!��R)��A�*�����P�CH���g�T�,�&c��{t0L/D�r�(����<$Ѱ\���.��i���Ɋ��&!�8\��+�J��]9�˔�M "�=�a+����ԗ�u�h�I������8J~�����i3V���ÀM�F��S��FuA�L�x06Q����p	r�J�-�����Q0�%ay]��U`�?~arxPV��'V>َ��,p2FI$�y��dt]�T҂�	���7��� �!��P?Y�~Hs�	�.�{�ﰊ�wy��?#��3��Kc��|s#��#�����N~{.9���
.�H5X�|�f������ ���j0�#"�O������ó��vo_�q��p!�EB���ߓ�**j^�Pi+�Rffx1��%���I����n^#��}˝��O��"���!HܧI��r"��_����W���Q!�PRS�SW�Exxۯ�6�P���|�2��*�V�8ސ��-?�|_̶��o���OC�b�H�Љ�O��ϓ�5K��e#�#��;��!�7Ϫ��h�����zK��k.�&��*��U̾0�d��gƓ�[���%�j�7q��R�����Ó3����L� R?/Vh��kf���jL�Ui��L"�n��~�v!�j���0�.��e�����q��A�U�4@a���{R�E��D�۩���M!'�$�1�9N=����YVZej>��±��3�("�����+�����p~ޱ�r�`a�D6wV�e�D�IN6b�%��+*�������!+�9���n��
��$4pOfkr�n�m�Ld�zQ��$��q.b&�o�Mv���Ѩ��,�^�������q
�r�I��a���i������y�cG�ŏLt��˧���R��*�!b�G���	$�کO�^�u�1��Q��8Zݫ*F�z�Gp5��C����*��W_d�hӪ�F��8<�Ir�p[wf�:o`9�RI��$V��g����<){��i"~(ґ������Z_�����-�l��SH���7��Q&c륲Ȣ�Ai;q���W���{��oqp�T�]	��Ym)%�o�ӿ[�ZO��TB8�9o
C�\��zk^�7����y�@����٥R���/�F��u/��#��NA�N
eٲI�/Y�����d�
��B3�
��'�}7��p�~"Ih�1%.3`+���D� ��]٫���BXF�;�,;�,�����R�/�;��".�6"��ڊ���b�L���?�^66c��|��$o8�ҳ����^8"83�����,����i�o�q؇ڔ��}�|Φ���.�z:�ɽ_A�S��B�+T:�3��E�����8�M�[h�AJ A0�����}5�664��΂���xMZ+�X~���sQP�g�u[�X�=T��aE��_μ@v�I�g��Xi�F��� �#V�����^���ҷRDF7{�z���AF��˕�2-z��au\z��ӽ�6�����=�<�.�}d�fk��)�*�-��;�N��1�9�g��m3:����wHz�mE������!����O��yYu�B��˰�HV�ab'��J���6�T�5<?�Xv�_�(ZY�.x��<N�k��G&IPV?A��2eZ?�*�L��h��5
�V������"��͞3��p�� c.k�{x�l�H[�~���|�GPLY�P/
�H�/����b�!|!��Ps,'UF_I|G��q,�r�Q�.ʕG�UU�7�����`��u��^$U���BP�������K��9��p��1�:a� �j�=�@*e�;�R��˓��5i(���l]e��9B�cqC�$[�vy#7�U:��V�mM�n�D�"�h����#���ez�����	���7{����J�«����N��cG3Z��=���8�ș�����c���Vt��D���3�?�c�qج��-���MS�t�T��~Z��I&����$2L8K��p�7*6:3��:9~�k�X��3�꽹�$\�2�X�����ߐ=������57]��W�S���U��������6C�Aq|?�5�`t{��hF��=���v�dL�!���(��.�gg���J> �[A0ؔs�^�	j�vژ�pBz�[P�_/9-\l�ܲ�X���y�E0��0��.Ż�����~��y�����.�1������,p��8\�w��4Q$�f�U۹{��|��O�)�$�<L�&��q��̔�ԊM��'�!Cd� �w��H/��� -��b�H#�Hd5t$�zi�����Pχg~��w��=����y�vT�<{�35�eR�e~
m�;�Yp3��;m((���;9��~I�ϵiEyWW�%1Y�GU��1����@y+�H�@��CJ	�ȝ�F��3l_ө���EZ!��?����/��9��-�#��l%T�!fJ?v~^D��3��.���+:t�	魩�(�}���zU��p!)-ͯ��2	��] oALЍ��o�S3V�%'"�]�D���H��Y�>5iϝ���F��
�H𡸭�H�^�s�h���1��Z��_4�mN2���7x���@�E��E嬨�Z��� ��0stj���I�1�͖��?$c�|��j�l�	�;�I;%�P#z��gs>�n�D@�<A�h��G�C��q�ᇥ���ux���)*hԈ��춇G@�Nl�b�cԻ��_�a!t"Z)��������O��'rץXW��#]�{ߌ8 @ߠՄ�-�mr�Z<��X�YP��\�U��bBZ#-bFf)\���AQEųmGq�ⶒ*��H��Z;r����� �٣��:���r�b������6(�>��A>1�4Pb�`o�y��\kV�V�G�T�w#���Q��B#P�x.��q�Z�c���-Ex!�l�F��\w���⬩�8h�і�(u�J?���P��OO�F�c�)���r�̩���Ó�Lߥ�G?×L��S|�:��Յ��&�!o��hZ�V�r)����P��H�̙Or���{�
�
��8eq�U��b�?w�����y�vj�%�g���^���}O���]KKD�,�sW�� �ׂ/���z����kok�x��I���SD��iA�<	qmY���֋!��\Q��225t������O��m��"%���)���.rv����Ƅ-��#��ڹt�@9�~X����y�N{��O�Q˒*� ���[hd�Ŋ�|��~V]w~�A�}sϳ�!��ׂKP ��yfb%��\Î�ŝ렆V@[-,j�R����uŧ���C������4��YX [&�����	�=��z�@5l�c1���z�FC�n(�����i����[q>4�ޥ���ċ򿭷��uƺ�tїg�Qt.��\L#��%��U��'�}�G�����;�x��/��ݚ7����M����I�%��jG�&��5�֋���wBQp %"-�at���*���ɳ봭9��8R����y8��CcE'��85�]�����#��=��Wl�ŔY�^���I����`6?�o�lg1�����EEF��z��m�6�C�%�������_��RV�����*-�oo���>�l/z{�5�x�P�7�����o�ɴ~�������c6��＼�F������V�hi��-uh�&��Q�ه;����k���$6mK?�3�-T����� F�PJg���(Ǭ�ލ��yҘ����U?!e~"�cY�Tmv��g��06�����t;�&RN�6C�s�6�Kfj�I�Rs���#ىuh��6��P1
����K]{m��S���,��C�V�rNq#�<�Z����o�n����+����J�^���G����j����,���DObiC� �6�TU!~<2���zd�¥H~<��m�ڀv	�����^���Q,�dc{���|2cy'�������ש�~퐻<9����eqQ�67�i�=,�`5��И\T��V��������L���n�h������W���x9WսY�2���c�<�ϘlB���+�p?ft��6�#�D�����Ű���ҌZ$j�o�@,���ؚ[f��*~��d�a�f�H>b˨'�M}�.r����P7&0bl��l3�y�]����8B��4�1���p�6	�$�<����	���r�rs����~s�вhv�Fd>�������֧֭��}���Q�����6e�@t~`����L(����ؒ��5���bL�n�[{kQ���lf�n��ym�rp�֎f���\;99���(��l^ʞ���;�:��蟇�]J 𵻅^�AҚj��9T���8\�3�����'1Kj��J��	���&]�͂FQW����+�#ke���)��ogV&�B��th��c^!�����+��j� qww����N�����Awww���!����߿��p`�7����U�z�p�.�ۜ��x7%+B����T�K�������+)��(���^����n�b�w+n��=wmw��8}����bY^��!�YbI�o��3�������P� ��V{�Jj�v ל)pJa�nGQ��>��R�d<����,b(K�o����ܮ]	)��٥���.b�~w3��3]o���m��O��=f�WI+*�/���r>���$���"��N�d�"7�;vV�uŗ�z���a�V��=$��P�^B�?��Z�A��>P�Z7�+�Lϙ�8�;{����;�8�$�'`?���Q�_>�)��T�6k|���"S�kF���,<��Ltnĥ��4([C!}$�--�Vsxk��r�%�o;��ۃ��3Վ�i�n�1��&��'P�1�F��L��yfc���-N",.m^%v!�p�$f��F�}���kO7�(�+��YA�������k���S�e������]�Hiii������W..�PT0� ⮩�f�M8��� ���d���8x���)� %ā]�_�~�ӖQ�yv�[�BV��V���	M�-���o�x�D����lxPlu�����@JS��n�DPz�++H_���̙�M|}˫k2�}�D%����)�#�7I"�s'�;NF��)!�'K�IX=�/IB��م�Ӛ���QĂź���T���>p����.��K��( ��=���pmm-���Wc��C'D`l���G[�JT����Lh��7��/?�.|,�W�pF��`_ �D�>o�����0�4��M���#��7��zj�{�޵4%�)tdki�]�>�
���Er�d��:Ҥ�y��[Q[7T=�I��<^H�c���YC��8#�����,������"'�<Pj�B|V�~�Z��؛ӑM����F��x�8b;����P6��ï4v��H�V�y��Pa�---����u	!O��P����5-���I6X����-��yvV��e�!�QN9\�@��i�*Y�!|�QJ-����_���[�X�@T�T�`g�,^F�
,z���%FL�{}�=�W:��{s�l�d�r�a�n��تL<Ƽh�������#��b�����0H?��n]0y��eMt�i����7ڧљ���Ȥ�L~�3D��',�ۡ��n�k
��P���?<�W�6��iI����[Z���pp`�HΤ"�*+������P:[_)�& ����rx��%��￪����o�k��o�uF��PLMM�ă��h��tf+.��!���c�=N_^�ir&�����EH%��B>h�5��I0t�sA�=�u��DB�cB�qm.�/h�oũ�7��K���SsR}�^ę�U�c�Ѳ��А�u����uБ�����7u�V�������0Q bZ or- ����I2r9u5ҥ��sf���ë�����c	
���Y=�/^?4���F��]������F?5���j�U�����'��������tE��1!�K��J=t����M�eԯt��< �ZU�V�:��^$B�sև��L�[��@G�|E�|���/i��}�Η��_���*��JuA8x�T����(nN�/��y�S3\jX$Z ����e��i HD�V��Aa#��K�R���즥T���j�I��cj��sd�y?�&F���IJX_�'v�wU�W<�[rj�,KPLFl�i�a[{��j`H� �0�D+�X��n<�ʽ���"�d��k�O]y9��:���9�ȱ��n�v���T�r��_�x��_�����
�p��t�ܬ�d��<P�OQ�P5ăA5^yՈ�:�!ۇ���j��;p����{T���t���B߱�A��)�s�lo��r��Te�F ���b,h����r��Jħ����zT����:�� t��X��i#���&38�:ː�	�n�Eɐ=lp"�L�� �"��)4��=�����
c� ���A�6��[�1��m�����z�ֽ�{����.w�L���I��k���I5� M��T�������K|>I���d�	o�J���圁�c%C�Kio����y���N�����zF�W��Ӽ �!ˊ���8��<k0���<`����Q��ǖ5鉫R�D]����_!�s��[�8Ȝ/;������	<e���2��N�Jt�:a��V�&��+4��D������S�p�L!�έ�Ǽ�Z�G�Q�q�b^�0<.��2F������8na.�ta}nN9�,rwB���2�)J��5�g��Ks��كU/
Es;�q�k�4",�����%/9��ӗ�&�d�8�b��t��V��ݥ(_���{�K�B������j�,mP3�@��b��- 7KeFFщ��
Z�v�Ŝ��ضJ������!.�3�ʿ�iyԢb`g5� ������J��_�o�$E��L�׼"�[z�OUj�n����߫Ϙ�t"��I����%��;�Y�@u��KG�SOG�1ăVfNKF�SF��Կ�pȍ��Bf��Ahtn%Q��9���D
��R�:��X�]n������`$zm���|g����ؾ�q�K�̄��({��@�iY0F�$
��=�Zi3�qE�,L7���|7z���zј�f���c�znIL��3\F*�Z���9!#Z<n:n��9�9&〪9s��/I0�g.x�NȤx����*0e�b ޺�ĖT8�L��\A�ʈ�(�g0�������FA�Q�a	ѫ	�F���y�e����k<���ۨs����@]��㳻hA��$û��fdk���~���,����+S�R�4�:���M��ú"z02�q<�k�v�ʑ�H���U����p����iLI��Vj7�;���cI�bs7|5�?��*j�\j�ײ�T:�j��\͌L4̇�Q�N\������/��k�`;1�����4 �G�B�g"f����.@AVhͥs���r�=���G�?ت2����S�x"$���h<$��Os|��nQ�{ �x��Kg5�b��D�ڬД��xJׇ�1"M�C�ʬ_��]c�T���`�V\ōy����*B���9+�dqW��KR<�i������r]x4Uw��k��}�FNb��%�qt:6|*��P�{�O�s|�LP,�� FƉQ�La�y�&U-��u���@���Ȅ���p�n^]G��&{VZ02J�%�)(0Qc�:fb�ķ���@�i7V���3�u��q1��\zؾn�Q{\�T��b�Ϣ?P��8�܈#�D����˿�W�����u�tu�S�B�i%D�l����P~�Kt	�iRF� D�1�-):0|� dpa�a��w�U]W,l!�<���
��F�H2��U.��,�r7u���.I�c���,�pV�"G�ee0)0��GA��Da�|����Ad�%����r�dɄ3��p#�#㇀&��
o��1��[^���U
�f���c0�)�L�A�ą�de�(�ŉ5�~�CG�Gxf�Z�#��r�D���ķ�F�S�N��jG>f$S�WF�TP����a�_W4I�*�׻j:�yA������`�j� t�$F�1�Z��ʣ��x�����8M���g�M)e�e�sHR�Jit��cR�� h@����Kz�u%��+���� !�����b >��H��(�`-\D�b0*�(yT��1&������a�����.c��7���v,_4�"�����߽�ĉ0)'d�h��_������H����R���~��=�+��H��T�	��4�~DZ���3�F�����뿘��z��H����{%0�1Za�p�t_OЇr�>g"�[�6�K.�*���+�FNl����q���k(5��F.�豮%�0'��f��Β���&�C����G��p9g�`5̨�gnFR�	��(���;U&}>G����1h�	����tp�b��!2��3�v�x���G��ߡN?�P�-|�ߙhK@;� ��33��<6V<Q�#�_Q	�8QX2�e��%ѝ/V� X>�:�+����o�6h�Nk�=F�YnFt�AKC�i�J����ލ&��Z����rRG�x0��*Ng�ܛk����� <M��P~M@��+�\q0j]�jG\A��=HDv9l����-�m��i;ziZ&GT)�;n.*g۝�ߓ4�ɐ�(���D���	��D��|�E�o�"���C�՜"��)��NF��|�q�|3Q{�(��=�q,X��\�f�s#S���}�MW�	]�:�zO��ޜ�Z�����A4$j�%u��wPh���U�������J?�'�*XPvH�Z�H�̱Mw���L�V�� �&��F��K�*Z�x�j*T�o_ݥ?������cO��
?(т�^6ph���5B�W8"~ȬI�'P�<o��ʱ~3M��)���؃ �1۠|5M #�n�r1��k0B�W(�x]�χJ�Z�͟��p�v0t������� �}��H�Zi�����=H��=>�( �tQ�lCX�W^�����L�d�gb]R%��i���}��O�d��Wa
;����Z&���1/^)��kBD$�N����Iq��gߐ�ˢ:�{�=M����&���%%�����4���9޶M�(8YZ�Zb;�|1�9hfv�G,}���4�<i�ѐ����m~]��M�g�oĕ!^}^e�%Q��$��z�!Ѽ�&G��,��H���F�
K��ϻ�)s��HO_H�3~��c��bj��̛`�]��	Vz|
B�����t%b��詫Q�������ҏZ�b����g6ܒ@�i�=�I<$u��X	��v�R�6��Y��
S����%�O�Jԋ�
��g�/��|��]�/�g\m�I�Rc؟�YJԋ�@��!�؍;�E~���i��L!ar����,��x�o�7�E8r���<6">]��_�BS��&�	6�w����Q��]e�E���Ѩ�E��������� �H��������m1<����ƺ[���Ӥe�g��	�� Z�d���$2
�J���Ot ��NCTj%��,g {P�ɤ�Xs���Y��A��\����Ru �`����˕��/cGI�tE�f�TE��A8:��*Q6�y+�|����P�j�q@�\n7���P�J.v"�k����v�R�p�D�Q&���hMoQ.��fQ9�X�M)rتt$S"�n2��$��եwmSm�Q-)�^G㾌nl��4X l6�ئ�l]=�����rbS*�S���)�#���8���-�x�qkS��~vFj��t��(�fl�v�6�y,�b:���f00�X�,�k�XLţş@<6 KE�&��6E��hOe��z݅�	��̟���<MF���T�V�y��)�%�5$�����u��Q�k�D�	o&�����.=�p ��@��PIϞ
E�i�P�U?�&��2��S�U ��!����<�� O�q �Te�wlᖽ�ܙ�״���>0�u��g=��ns��BP��D�OB��|����<��*�@'��݉f"�A��t���+\�6��뤦LCm]M!ߐ(�35���2,�MT�������VL��?3������S�YI �G�_>�f�76� j�K�� �3�DW�L+a���C�q��,=$����_߻Q�Veqb"��k������n@o<��7e�$f���~�'��I�tN�	$��D���޾没��}r`��&�1tR($q����-*�����0(�G㏃�d�Q?$\���7X5Y���؇��fm!L�8	~�\��9V��Da~f�� L����ig�s����=���x� �84x8R��.�*�O'�OP��_M��HK���^u��x���x���L��X��1ߥϚ��$ܻ��wާ�ʧU�[]�T̎��j�G�u�z
�E��3v���9igeW����5����z=��������n$�X��N��8d�kqOqH�����m%�|,{F�������'�c���[�)n�]�Wm�Z·� FN!-_���X2�|pdCu�ob^��}�RfDy�>j� �JX5�\����*Q�Z��?��"�|��^ �:w�~�~�z�s�|D'Gf<剜i�����z�6�y[����6�"tw��p*�D8����y;E{��~'��ZC��̮Y׍�=C��U��ˢe'닮��ʯ����"��A���$� ��{~D��	Xr�8�L�\`�S�̎�c�؊�Gg��<̊����P� flL�jʹ���*��Oµa��+OȈ��T>=�±S���Ny�:��[��X����~�yC7><��{�h���:�2��26웈�Yk�x�W���l��j���N#v���=bܾ_1��wR���۟�S\k���||L��o��I���v�/���j�{ ����z>�,���D ���e'�v�G\8`k+�(�P��'��h0�W�+̤�j�*�qêSu�h�cu13*�D:�N'Z��!���A��E`���O�5C%���Ꟙ�{�z���Y&���P����?���wF=�o[n��7Y�p5ԓ�U���`��b�_F�U[�`��3ǩ<M��f8��](��c2r@t �0����.N��X_��_�Î�*����Nn��ȇX�ݜ��Y�������&�P�S��u;���s�I�k ,8ks)j���������}� i�~#o�g��~�4��]{=�*�Ki� �!8����=�1b��}�1Sg�2U+P2��L�˿C�5��`vu��� Zv8"T[�r%qW˝�D5L���D'�4�~6�,<T%�\D^^�h��o�1��#)w&�*jl#}%�����rp�XA������O^>�����y��ŤL�e�B���#}����2�=�}<��eḦp����A�Їf?\թC��0���4��3�-zN�o�Xy���rw��e��D�нM�#w����{m���_%�I��%���j5�}��)�9���6abT���vD'�i%A��0��k%}�wT��Ɗ͉���W� ���)dF������4�t��� W�0�=�Jj�\�,-G�Կ�Z	~�2�Q���P�P�iX$̧5�E$�8�b�R��1�7eh\r�+�!g���}�8�429x\˦�x[~�E��I�ؾ�g��8��`�������ha^7bFvqI��;:�0���N�lޱ^�o��?Еh(R��L��ȫ35C�t{�����I��+I�0zu9qII�²�-�e��fh1��H��`֩�d,�����_m��((ŵ�|p��ߙǧ��� ����Vx���[�����	[��b�������+W��ܨba)��A[�^�۸8�Z�"�������Xm��*B}�3Rb���y��z!N�B����%�)ma$��Cp���8g�\��(����'Vk���R	��k��R�y|��#(�$j4�Z�_�N�9)}}�;�+�#;��y(�Z�7`�%~�m�4y�Q�ɳ:K��\(��ݳ��!�H�6�}�ǚ��X`����.�G��1����׻ƒM��	��0!5?Tt$/7�eև2ɋ+jTd&&�y�ާ���5�gw�h{`�݅�\m�l@�T�:����Z�U�HIea���3;�M"����tеƏՌkQ��L�0*��1�6�"+q5H,�	f��ě��:7h��iE��η4;'���\���C`m<���T��%35gx�h�B<�d�P�i�lm�\�y�� KI��Et咿P�"A���l�2�t�����im9�J�`��6�߈y'_ڹS0@�-���7QRhԻP�\^د^�v�f"�>�a$u��-�	�[�[9G=���Z�=a��Ɏ���L�2���C�ZX�G�`�	���@�1���Y�K���S���������t�.���2�8FM��N��g�#�5^.��ِH���S0�*�ϯD��N�H2��ޯ&y����q��z�]%���򢍮�M<�Se����YJ
�;���
���V���g�k�1���_w9o#����߶"�>�/Mt��$�	q��F�|`�W<Y���s�34\��7���6��]���W�Xъ������HH�^�*5��C�ܭ�2���	iB~7m��N�Y�$��E��j��so�P"j܇�K�Z��ԩ���̣�`3gy�ܶK��� �� �ъ�6��g+0���o���t���'> 7�c��Su�����:��CƯ�������_�}V_���Hv�Db�䇪�lu9+�lXN>ZyE"Q�|�$6P��HBl� .���bwN�Xj�'	}���Fo>�]�:�/1qM�Bc�1=AX����l�~��
��N��wu��e�b�ԏ"e�}��n�,�5�� n��b���nwt*�(2���e��/ԅ�
�f��)�i�;�{�60�·��[+��?<6F?���o�~�ɫw2���޵�A�)KA���e��S��_R.#p��6���` �'?Iۦ}�.3�'�;!�"i��_��;�/fq����9E'ey�d�Fr��!�e�S_�D��@�����zW�ER�{>�).)u���u�B�*��w�������[?�����6;ﾛ	�o�����&s��>I��(�M��B��A��~M<D�↦�bq�W$�N�������<�j��M?��,�m����|\��G�OV'ey�[v&�p!$�r8��5�0g�����䣫�����L�P��cl��nv�;���}B��p'h5��C���ˊ@���R�j��O�|4���Z��xL��xx����^�t���.�`3Z��IȦ�.rsRI(
σQ���ri��;����1KfH5�uFEB2�̠w#:4xg����Y|��fJ'�j����&�h�����e�.T���D�.2�x���a�u�%q������fH���D�G��\�'�#�� ���+�+׻���_v-B�Eļ����k�[]v_���9���-��m�*Óf�׳�%��K��Z��ݰoy&�N S�n2g���<R�/4�]['��v:�q#`�?��L�*؎<	����V?hs�4%z{��t���}����eQ����)�;O�>�zbR[O+Ҫi��3=�9z�u?J��d-�AR�W+�,<ؖ����9Ӱ'���Q�Y��9�b��?Y���
��	�'��Đy��Y�v}�X��',b��o�x��p]��	�O��X�ҟQZ-y����<ʵycxU�T(@A�0h)�����0�@yh-[����%D3�V�r���3HP���S��ŷE��#��FtϾ�;!L*,��m&U�i;� +�B<� /��H?�l�`�Y�K����p��8�=���v�Z
�b��mt�&��O��Y���r���]?�1��o�w���l��ؐp����L��V`��d��%餓�&�������T?.$�z�F0C��e�by��p��$���F_�X%ϙ�����������	�?5���ml�z�������xU��~�������ȼ��u����g�����ޥ
�,f����jsU"o}�LGٓ}�^�X�P�x���hM�0�4B �cS1��o�s���ݐ��sd%��Yzl�ģ���9�*`�kj�kNU9<]	�u}��o��B=�+>z�Fr��_l0�v� ,�y]�?�Ѷ�wm��-!쌡Y��[����3��������B���t3�K7���#�� !-ºK!�#8�s�*���Jp�ۗ��dO�a[��[���" ������ǄşC�yQ
��<#������X�����I9-�ܘ+��Ȇ.Wz������D��H�N�7HZDW-QK0�.̊O>ϻ���Pt�Ȑ��B\6z�՘�D|po	�X�'J)Ϭ��1�svTӣV腀~��K���S�NB�83q�zJ�ז��گ�á��r�o�Q���hͧ�|&��0@��S�j���|�{�\'���Y� _9�B�O�P����+���[Ԟ��gš�u��BT}_� �J��A���O�X/��)�p
X��% ݂�	�� �B��
ε�8�s�gF�I"�S�j�w��j�q��?�E�(7kOO�1�m��`m-���K��<=�ѣ�t,��8��?n�zQ�Zʙq�ˌx��A��z���=�E�H� r�[�(t�7��V��K�M_��P��(��ة ��c���x����$L!�D�j/������#��'!킣]�]R0��^9H�*l���ӽ(�F%��'�:��֭�Rf�C�r���4@F�S�_>>��BtU��t�s�Dwe�ި%�������T�!	�d�3sm	���(z�?�G���R����z?X>��0E����6��7����C[�;0��u�����=����Pb2�����1e;> x���p՝��Ƚ1f�q%��p����'ȫ��b'�J��	�>F$/�Fm���P�ˑq�_����HQ�A�i��V.�]�-?�*�r���Q5�����a���c�K v��^��~DS#;�/��(��~�����Ϝ���&e������\��R���݋����^�z����jOvS�F�]h��-a*/��T�J�eFc
N���~/ˑ~�Z%�s1�L��/(R�í���н��Q\���ҝ�u�uT��ܷ P�;1�=|��5�U�L2b��{L��$������!.9���!+(���Z�R�� N�-��S�`�[���^N�;L,8S�\X��s��0�JG#(t��ޜ��ޗ0C��O��$<���\]5u!��i��=)%��L�͹�:��z�t6w(lW�b�Yn{52�L�f�4����
�.�8�ղ;��g �:f�d���r�m�o�V�ݜ�'�	����:���6_�\i
�����b]p�~
 ���;j��,.�������f�S��b�\u��:����Nl}��[��tE��jČ�{/�f8��)b��EA&���@ļT6�axXퟔ6� aRvgjtV�H&�+�K3o;!��Nkz�1����Tk����oN�P����7���uIl�,����̮�i8{z��K�'�U��y�/����,|E7z������zp"�?��z�U���k���|֞wBp�23y��� ɶF�2�(x�N�[�@B��LM�-�K����4!2�����e�h�W����G{پ2�ha\kĎ_T�Mힻ���d�X�7t$�́�__�c�rÚ��P����ƀ7��Yϓ��y�0|�> ��a -�s_��ȭ��b]݂S葩��|81B��C�5����֤:>�K��,GR;>�6/d'�E���(�|�T���^7���{:+����L}�i�.���ʟ̸VF����{�"��v	��_]�z�~K��Z�){ի+Q��'A||���l�/�2�D�9��'H�;��;���`4q������p.���$:V�ʫ.�� ԝ=�pei����i3�m�L���JHAǞ��K~�ֻ� �����,��T4OD�N"ʹ*V���5q��/z2�+�����TO��D����}F
6�I���/������l��p�D�4W�Xѳw�{V0t�|�E3 ��ٺ��]�D�<��g7�I�(V2|�z�[���m���M� FӼ�д\�]�}%5�N��ams����֓��?����r�E���k�#x^�<�5����
ѧ�4�"8��^u�l�����4]H�$.��Y�?�ŌUNT�r�IEq����Y���}�n k�<�����^�W	�w��ED"x��-��ʬ�����K���ZV1oj�0=;�{�����Qz�͚R�c%�ps��VX��5��L�W��L�i��������D�rP�R�3��&��]&|������b�HQML�0#Em�p�zԩ)���Д&m�Ek��B�)V$Sv|7��iҸ԰]i٨�aI���p�D�&0J;��>�P�ɂ?wo`�-��?��|���?O>��R�y���>#���L|�Q�D+���ei���.^$t{��&.S�֛b�;A��`��#YƷc���A\�8���7njp`O��ֻ���9�H�]�O-*ϯ�a�Ajj�#b��������@i�۰R�`�Ǫ�i��˭Xy��
��@D禉c�1C�ޘ�m�+��[� �ǫ���CTw�x?���i�AK�~*��02�3����T�Ԍf͡}��tz]&��ސ �h�n�}�J=8�;-mF& Rc���B�H@<�1�,uGS�O�c�E� �6��Ƌ�tN4��{�.Q``��z�iP�Tfjڮg��JKd�ع���u^.�t;�y2����4��e�A�u\/������3a3a@�I�b��V��Q�2�=�{���������f�>����`��[~s%�[�,�//0���V��~X�8X�v"|�a�*ணf��_��6�	Z�HZdqrO�?�n�-�I�w��6�/u��!�6�j��е�	�J{ �q=-�L�B��t�W��;n#��f�y�rÿ���ĿR�T��v�ۮm��O��=)�R�PN^�������f����z-��nC���B^��0���#����Ķ	e������שW�j�e�uX$�[�s�ß�S'��g� ����<��02e߇_��/��YA�HA���b�
� ��O+=����LȞ��-52`�T,n٭f�_tb$��!���}~�����l�LQ���9y��݆fDp� �]:?��}M���Ǒ`1�^[5���\P�bu��Aч��A,�s��7�#N�7G���52|7��<=}S��i4(�D�K]F�\����9�=���YyT�<~)��ft�>�ּ�,0J��y�Zp���@��.��ΉgS��R���:&��C��+���`���"d��*��d`C�'�]\��}`P`���� ��*NA��hj����E܊���ٓ���@
�nm��J��%s�Au&�%WD��3��Z������BB�{��V|H���i[8z�k�	#���w}��]ZW�b��G:�Bݭ�R%��������JB2֑P��~E���P9������\�d�������E�b��)���g;Wq2���6�=$-5��w+^O��R�%�Oi�^��$ϕF�y����:D?Vi@h�bi��o�P"���t��� �n��=9�{�d6fZ������i�o}cԦZ��~@��\��v�����#�%,��x��Ɵ�����9S�O����`�aV�O�tBw���y��Ƞ(q��"����"O"�?�[�p�p�RF��gC3`f��#��F,O�K%4pp�>��y1�)8��
����+��o���غ���8Ko�8V����}�r �J��L��,>3W��Fd�K�E��Mf�Q�R���١��nt���E�"p:(�-9�Rb�M��h,qU�$F����_����%��"��[ӽ�����4k�ղ��%g4Ӓ�tp�Dj�rs��	�aT��T��'4m1����`�+�48c<?���2��`f4#B��kJwhnw�X�[M�!�fsԃv9�k	�ԂA���EV���[=�:���Aiɨ�TdA�N*b!�~
�:�Zu�H�b@���=dZ�EJJ��YDƀ������ᚷ�s��!�g���[w,�f�D*����qU*E7�cAi�����4�=���������Ax��uw�4 &�^�'�Q��]Niu�ƈd\��NS��ɀfo��*��?Z�T��]�r8�OlW�f��̬�_�ޜ7�fP�c��ҧ|^5�?Z��(ˇe`	Nu}�cp�`A�V���7v�ӑ��yi.r��b�\9n'�AV�j�-�\1�n\���J�"�
e��?�����ÿ��#S�)��kdWb"�c�i1��d܄E����.r06��feܯR��V�ǯ�k�����W֥��L�î�[j`����#˘��HJ�����������=!�'��w��5ր� d��׹����U-�&M��\��=P\_�9zijf�-�{��U���(�Ug�mX�v�s�)���q!u��	�l�p�߳uW�8��� J9��ND{I�=���BhJh%�j�m2{�~\�5(rzӎ���PfG�њ/�W{��/@��0$��q�!��n�͞5���CyƏI�������na֤��P��_N`C����=�U01Ћھٮ���ô
��f$�:��P�k��I��Vg��7���E�dQ0����[)�y�z9�A�v�$�j�w���Ǉ�&r�+#����V�G?����'�B)���OQq:�LBr�E}������`K`��1��z<��HPe#����Պ���Qr��g���8x�x�[�Y�4�d�E�`��.���L�c�����ّQ�d7�jN�CL�	)����e������kM#�^@���J,��K���o0�e����wEy ����}�q�������iI�|��h�������2�(�����6O{-@T3q����7��۷yu#~��j�,`4�Y;�m	�cϷ�v�Bm��8���%��%�A���qo������B�@P����vs�B���h.��@�ˎ3�=`)Ӄ�;x�lk��QɅ�OK��I�/����n^L�����ӵ(�ʝ�b�V�*(6n�q��bb"�W08�ޙ�>n�zj��N62����f0_��A���UE���r��W?��y��v��{&}�`b�Y���b.���,����9p�(� q��~�jdl����o�b��BX�1�OE����Y��v���?��Kٷ��P�b��&(&U=��)u_�_��6h�]���4ႀܾ�U�:$�G{���GYNK�q�j��CP�����X��!�k�_�p��"&�N�*����9�n�#�G nq@=��J+x^�$�<8����SD�x�ޝ��@E���0��e͞�v�ev�<�i��ܫ��|��kb��T���xn���^9�Z�����7󀨟D���d�w�Z���\H�US�4곁�!JbC��[z��^7o�;�{�旞O����}��|�<���3Ç��a�P��fo��a1���c��6ҹ޿#�C�,Ȫp���A���h��.��J'G��)B�S
<\nj�¹��k%j�.s��4��5�}�,Ȝ�B���t�F��"?�0�vW?Nf_I�?��m	:�7aU�z)����thI���\7�޾�T��׋��
?��V7�$�z����ɭ�觊�����
}�S������4P�H��+�o^-w��D�!�Q��V��Pߺ�>@�⺖����s�ϰ�e�g�%��'����=�j�ζg��fďsˉzW Y*��1�>$f Dx��{�q᎘�
s�FKk��a�B�F�aO	�G���n���F��>���0gEx\�;�����]���i�[6ˠK�4��8���;H"���~���MP�%OH����M�Cf��o� ��s6��yq&�j�T歫[��^��A�3�KSS�^׆�HgӨ�4ԃl<���y�Gfmχ�=H���&� ��2j���A�X���z+(��͇<�èb�)x=bth��$R]��# io����m*3I����0�NPz�>=��4D{��3���(g��`���!�Q'G��5�W�_��|��	%Q�#���5�n��D��R㮪�t��-E�W��?�M7�C3> �Bn�
Oy�U\�9�ָ�L�Ń�jm�b��)D��.LT���Ί�=G�A!��'f�#�O^��Ԥ������7zҸ����+Ϻ���r��-�Y�"zk�z}>�5�a��3����뤔F/B8*��!�2�H��u�@�iOd6��Տ��߾�MN9
�+?�etJ��4���;��w�/�J$b|�׏:m�C���MyX+_�鮳�-�B��7w��	�J`��\���uw�Q��(�-߷�ک�+n���G�]Q�� �����
�9Tɑ���YY�^kKѸ!��i������6�'R~�
�Vb~��:��fAD �<z|(�z����T�	-���๦��Q��}L�of���T��fmgm��b���3�G�`8.,�=��ż���쳿� ��rŤS]��D&}>�϶�ܗk�R�k���Ee�{�,���Wv����[�6��U��:��wu.ln̯��-�>f�8���^�ػ9z��pJ��Sz��ݍ� ��	<�.����'�Q�����j�E�J�v&ɥmw�A�ef(0FB!�ڜ������u�m��mz��Dڴ)�3�������~s6(��b�*Zp�,�v�3� 6�``���$`���Da�d�2>z��?K�������dI�e�\!&�vʵ~<���3\Àh��t����)���oO��*⎬nO��z}���$��=�]�z8�OU��)�Nأus�!��
:	�=8���u����)����\��`��<��1��r��4R��Z�{����W ��4�^ �������!������	��w�<��v�|�{�
�����鞖sfzz�	�|w�mw�.��wZ=6�� �ջ��h�<r�x�D<n�͸��^�����\����=C&�vs�rȲ�#�[��߫�X�����u�.X�a}<�h(�/�	+%�q��F�֖1�U����	ފ��!T�\I����.`'D�ڶV�s�3��y��i!*���DL�B�#շy��������1d�M/�$�4�8l�{��&O�f�RR��{�z��wf����'�n��k�����������{j�9їӎZI}�S�˳[M������q5E5K�:�A
��sdwǪ_ie%+�W��0�5�"F*믖��և�H���s����_��-�8ǜ�~��`c+@��7��x������B���Z�8�m���j	�wv�q�!�� ���æY����|�1@dc���$�G��t�B�{PCSPɏw���4�BJ��C��җw��r�Ը>�5F�㺫V^>�G�6lY�l��@M�?D��kえ���>:�/I���Y����pp�K&�����w���0̍[We밚��:𮦗���.Α�\�v�� �TZnY �#�]�&eL����H�A���x�x�y��N[��h'�E��V�Zb���-D����|���x��	���\I:Ǚ3��SC��h]u�%�^3�n�u����#A�Y-G¯�s�����Z݁�����5�ߔ C7���$�~�C��!`�42�o<�!�Dvmr�dXP���y+���:��O��RT�Џ��hh5��x�VeKh!߶�o8Hi�Aꕘ�n��.�qfK��K��^��d]�Jt���`;��AO_9�e7M�4�s�Q@&�׽�L���7^��1J����:����%8^ RS��������{a/������W~����#��6���&M���mY۽|ޓF��I��E8���^�e�e���#x����ߴ]}ᐩ��
��#ף�������N�x���0��C�o���!A�M
�m ���]����>u�?:��zD��q�� ��֯]$
�������������ý/�P#�0֜�l���yno��q�8�GE�E1bE���K�D�5u^؈����9I.����P�D�����A�}:�Q�<~��8��l���k����k��J�if6*�Y3���>H�JZL�#kc�������R�F8�0��$]]]u˧@��i~��=w��x2�̃{�K��wM�9�^m�����.��]�y�/犞"}�̍�v4)�"
��.S5�˔O-�&ժ0ҥ5%o4	��9V�CYhw��KC>�Ee�gc΢5N[}���=q,Z�z`"��h:�
�J�ݽ�ܽ&8���:�`#~>ݎ>RQ^�C�A�ʿ��ڬ���5�o�E���fg^caipL�:�7'�Vwvv
h���n9�ӕ������<�~y��4>az
0S�pRo���(�/)�b����m��I�0�L����5T+H��z�>VĚ�$-��kXdו��!rm�T9bZ�������? �{S����+�l}� �tP��Aj�d$�sa̕�&5Q�3�&鶵��3b��|�죘�jS]�7���9eH�,t_��ٷ�J͛[r�QD�����C�lXp(�w񉉉����;��zY���!?��OQn�A%�
��YY��3���dd'�F�괫eddP}	��f�����Dx�C�l_�޴[��b_�2�@�3+A���YCz�?�X�.k�G�?&Y��`D�؟�L���+nٱ*J]�����q��١B6s�/MT�Q]�I��*D��"|e)��%�#�r�WQ;rC-,[؊j��a�<7wwwS�Y�OxH�E��E�$]D�?�c�>L��V��oʗsF��L���zvnH�W�"r���@���<lדwu��/:�����J�ێ	�q����*�^ ��;�+8��/k�̓�j��Rr�]V�$z?��qD�uB)�<?�d� �^SZ��A	'Dnjl݃�ˋJln+"Ȑ+�4c�P6[*#�kf[�q��j��9ǽ�#�$�N��0�*��vP��x�6AH� 9K�	�ώd��xˀ�'�O��,�Hn�~�p:�9dn)7����5��_�2>i����\�d������<����o�7��9@�y���f�T�<VS�8�By�rP��d��ረ�o�UPQ3��B�a�0���͔+�p�ڎ<��+i��zA�YdA-�-ftH���&�*O���T�˖�7�d��O��GJ]��5wx�ЮI�.}�B��Wuy�^81o7|LT��D��ϼ�l�^'ދK�d�`��X�� ��)cy�,��"f��IL�֥�xgAo+�2Ej����[}K�3����T,���W��T���c届�vc(�	���(�햙MS�K9�廻@���~.2c)�����=K>t�>`�q'�d��O���.C��H*OeZ9�>Am�}�y�{X�"Չ�������uC�廂wN*m�JN8@~��X��bE�$�����a�%�
%[t�0 �(@�ӫ�5�U@7�
T�|z_��/��rY�1	1�kq���}�7����������R������ɘ�t3#���٢���ྍ��MT��:�^�a�:�2��"�ܞWu�7��/�3/;h��a��|9�טL��k�$��ׄ�j�R��G��c�~
v��L�Y�t�p�Ƹ�E�۷<} 9��{-���]�L�A���N�d��++�`g�h���X��#�t쵼��du�.P�� �xb�`�S��H�%;�&H�<,��Tds~G�#D�bF��v��ho�R��}�@m''��'��?<� �#�+X%Xg��r�(?;���ճr���jw�V�²O�q�w�MTE˂?UG�(�"h�.��[�����;�N0!}�J�G�,1/��^AbІ���˿�8���a��e�FY�3���;���܃���J��s\�����v|{����n�(-�1x/��V7�l���
��?��@��}��7�����M]Zk�[I{���x/��KvT_s�	���O�1>S��9�*=Ls��>Ϟ��[�EO���_(�v���#�2q�/��}Eh���Po�N��ozJ�+�(|~?%���'�c���~�g�V�o�9�:���#w���O����-�"��sB�5M�j����G�b��w�`"L����[ȶ]5���.Zs�'F���ԅA"5�zUhuϧ��;ᬿեA�9`�ć	-�Ԇ�l��1���.�5�Րy����삭��������L�B )N�7���Wo.e��^���)'=�h�D�k4��s»�c.h-�����ףc���h�H�l�#
��
�~=���1ӈ�_��-N.�zD�7��It����t�cQ�
 �$!eE���:��B��bcʈ�nM�(n �$
��uZ���l^;`�2�{�wez;`>�����]�F~+��_�*E�r^�xF/���\;lx�N�G7�7���I�ȸ���%�U����C��pe��KC��G��3��?
L6�#=�ʶ!������:bh�?��F�	0?gZ>{ĵ�ckK�g�c]",�l~ $��Y�wl�ԾX<�vh߮��5���dh��0A���MS�L\I���׵?R ��&-9@���3�Ƕ5aXvN3՚P?���~/�2/�]���̟�މ��.ӴQ?�v/���H��/GyԌ�r>��VjZ�%��}&����y���X�-|�x���I~��,��mЕI���g6xHxq�a�<Ȋe��n+������1^[�떵���b[k��a #d�����3ɪ�d��X�+灟�,��]�GO�j���\��/8O:���Ž��l��$�r�_)�:����A��>����>oTOM3�Ŷճ`�Xc^m�Uk0=۽9=[)I���w2��a\�O�C?�Cn##��_��c �U�V��Ύ��E�ыv^͏�F��0hq�}��
q�:>��:��,��L��(�^u�[�P�(B`�GW�"��D�7�v�f8�#$F����h��߶	�
jT+
�i����<;V�t�r��ʵ&��y��+��R�|�3����m�3��k6���L�%�C��������T����3&�}��A �7�N�;�8�hԓ�i�P=K��S���?�4����Lc���'D�V���N=���~��4e[�xV�J	2�܄�`�n� ���e�k�?�?sj��.].^k��tğ�v `A�?N=I*��k"��(�1k�SE��R�B�d��9�\d����@�8	�-��q4��	'<m_|c���Z��|�}�}3\�X������ D�i@��a�W'ǚ�od�����A��ALB31+�Is�(�uׂ���CX����� q�GD�bע!j��G�z�J�|gΞ#�T,���'���u6)�EQ!��VB�Y�ߋĪg�O�KQ:!�X15���(oY��FՓ h>�9���]zy�sSɴ�Y�37� `z	�X�)EX͛^ZLN�\Wt�lV��6�}�/:��c���I�w�����:2nL�èȸi��ʷ6A��%����i��e���Y��_���[�u,�'�M�Qr���V�)Wh0�nk�6���&�׋#ߘX�H��жY|��`hB*��j�RFp����d�Y�Ż�"���'����Hg,�7�-��N%yn�S "ol���{o�F�8b]���j=�N��Մ(���[!��|?p�F����Cl�b��@��NBX��B��=M�.A$@�'Y��ķ#O�(�8F��le��`k@�G�V�:?BR|��.�5>����Ӯ�`�;˲c�&?留8|���n�=�k;�Y�=���`Iаk}ۊ����9x)q���_���$��rP�TU�H�/��RO���~đ�z8	� aӁue�ܡA_�r&�g�J��ܣ����"1
LU<�Sۉ�5��˶��,j� ��8�<��{S����Z��Sκ,(!P��兮��b
�FV���Q#� �
,�W�8������v���(����_�������x����p���Z����"��[e�?,��}����_�9�FM� �2�>�T @�1��a�Ι�=�π���(��@��8��	#��A��P�p�|(�����sA��|��S�� .2��OV�s����P���
�>�P1W]����?Γ���l���U����cX�U�C���J%6L��3���a�f}W���;�&�`:��]�eYX��ri%i��>;m�8��vM�T�����2<�����<�暿���3c����M��H�<��@�&�}�\�ĭI8N�����D>�A��S��PA���I\���6m
s�gO;���z�h?>�KCJ^���\w�L=���\����Q�{��؟f�t�;� ��(���\��~k} �kM��ٸsQЖ������p7�*��9J�y��[������
P���Qf��Q>��ki��R��1�h�d���"Ku4�[�5����G ���Mc��ŋ1^�x�&7��,�DwNFF�y+_Hf�%Ƣ��[��q�j�����V-�Y��;�1'ry�?6�x�����&�Wҩ�"#�Ĝ���
�T�U�Ek��ï�'�������ul�_G������D�0ṕkD7]����_������3�Y#x���Ċ��d_������*���!�X�_���aZ<�8�Y����9&V�9�Kz����VW�O���z�kj��ϿԂ���m$�޺?D,����f�{�uۜh�P�}ݼ�╨N��>�RWjK�n^i�w�YW�H�'�	�\��i��"4���`����N&�e*A��B� 2'%�L���:��_�����s����1)�+�_~�nl5��|D�7�^�E��p�4]W�`EGm���eԑ�{�f��Wt�f?!{��>ߗPi��h��q��fX��v��v��j��e�)�w@��S�O~p��m�b$�+�i�>��%. �@�2Ղ�=���A���v�vK�"��&��Z���$�2�:ؘ�*ĬK-��Q��[7�#N���>���Q.4��q��]��ޢ�!�����Kf�l��p�o��0�,�� �E��v��/��}%�Vޏ�ȃ[Q��_��PUb?�s�g�\���e��.$�?BX�1?�m�|]"�3!�R0�TR��K�iBC�eHX_f_j!�!�J�l`��8���L����Gs���qc�oxQ֬�N��\�y���Nx�j�`��r+p�fj�t��H��$�zPGA�T�8��;���Z�B���}㤬3	K�n�#�ݮ�X�l�MC&��������H	�����}�+q/�Hx���-q���Ce<+�X��2�����n�&Ѣ6G��2�5�ח7k�9��C�ͩ����ɐ��/����*��Yh�۽�o4Kh�"1B���7�LGp?���z?o6���ح�И���q���F�dxm���`3��q�Z�R�:����"����~{Du�[#�P�#2?{�_�*��AnѶMxS�H"�Z�B��C�&�?��S�b5�D���>���WQW�[uLXiC�������<Ն-O	$��/F�՟P|�kA��e
Ҹ�M��]����x橆b�T��C���021:���-�����Ao2jc�
�`bR~`X��+N�N���H|*�@�o�ݜw�:2:�vlV��d��l�k�@=!f�G26I�QX�/Jra�����{6�4QF���^�����G>W"G0zs�qn|�t�C"�/"�1ˁ�`6y��6�����.,��[#�Z��D�����>��5UQ�ذ��-e���l[+S^�|���A\bLπ�P����S�O�5��Rrz�_6's?���jAp~�é���cC��7Y�mCU
�Gd|٬�/~O��ي�D��aˋ����CH����J=������W5�E�f8����n�ѱ������)���ֲ�w��*�A��'qQ�w�����R�x�h��#?�~�7n�����ٺn
4=&(�̓T��O�!NnRh�ciƀ��X��ÃKP�h��Ԃ�Ǆ��"�<A-�DФ���g1���%b�1D��i�����b�[���)~ݸ��	 ��o���R%��اv��?��s�����]dJ���g0�y�/�>�R�&'���c]�+���fx��j�����2�pq��q��%贪}Ra��H�ӿ���S/��[#j1'N���`Ǿ�:<L{8

�>$�����fzW�p�:x����8��\"�Xbo�%E�/�qz)�-[�Gp����6����FeR�ì����Z����'�YK\1��n
�����͜"|���p�p�=˫��~�Xz}Q&�	�m�dx��hL}zq��3{��빞:fPy��h�U��y�ӛ�i��W�!�b<�.{J�Uٜo'��(ة@��)�(�i�i)Χ�z)�zb�3�5��D=1����n��>�/��j�����f����M"Rg����	��Fi���d� � ��L�����SM%�61a���e��]�%=�ɱU����?!��Z_N.P6~=�u��^�o�X�U��%����M�k~�/K��@����r�S�+�����g�v.�z?bQ���q��u�f���b��a�����ݽ��xi�n��Z4�Rmw��.���X��o�ˢ�kM~�_�9+����o;%i�f�Gx���x����*��酢��	b�v�s��k�[���9uگ�v�[���&"��}>�+�?��bV�cE��ψ8��ao�D�szl�V�T�:�k��o-%Ġ�1I��rc�����آ��bKaM�Ye�R\�kM��u9��1+6������p����~ar�b��U3�=�~�䓬�esΝ��{{w����T�Ǧϰ�}EJ�b���'�[Q�σ[ҵ��M�4�l��߶9��	֪6�p�x/.3g� ���_2k߸��o�k;A��P�C;+����KOn���'/���mcN�T���4��t���!'L�L��6�R>�E*w��s%�|�7��[v���{J��_{�XX,����f6]��G��o���Y�m��5i�D��LG�i�&6	`X�	�B.����]��y���)�xz��ܶ־���rͬ�7w�M�'f|�Bz&ȹ�(F��¾�)6������E�ej�J�����g�������;b}a B��:��\���?�ɼK�&XoBj�g���C��]P���H�G����ǁK6U$�\�
	/�����3���a|m��B�Z�]��:����c&&�X�+��NOd澇.t?�u�R�<����j)PH�Tϲ�$��a��t��<��� ˿�d�� $ZM J(*[�
�9H�Ge���@J�M�Fm�X}k��=x��k�����F�'�cg
�1yR
�����"W6qg�� ��a��.�T1s2x�����A;�'��h�C��ɬԴm�*�B� �2C;��ѶL]�Ƿ�!����X��C����d->~G1�F���/�@�����}�Ot�����dj�1:��@�4�X���Չ��{bJR�D=�	��Ʊs�C�+��׵d~���<u@\ө�q:��s�xn�0���^g bs��}�d)�,X�t}����o0�����k1�W��k�[�6��0�V|^����7��2�����l�_�F�]�/0B<Zǜ�S�/ �!��5�`q����o#m��c���-^�j�r��-3<� �����U��88��r����ڱ�m�n���ffOA{�Ԅ���p�>������@p�S�X�T�&�*	�vZ�&&ވ�3y�4<���[f�eW��������&����^����X����d��;ʰ�� ;ݠ���� ��c�����;���rL_�G����6& p��:S�d�_��<��e�MH�~<f6~Q`����f'�ʳ��Cý
����4e��aT�v��*i�p���NB��ޠ��@N����h)�!s5�:�1���*o��i�%���uS��W`ʨՊ������j�G ��sF�I����we�$��d�!�Z4�G �=��HB�+\<�진f�Ob�����y�@\pMr��0ˢ*�#A\�#�^�3�D<�pkY�b����PW|l�=� @e)�~���qG�;��m�'��p��_��ݧ�����gfwd�Ε")��yj/z�l�k�,ܕhň���=�5���C�2m_K"f�ըR�f\��<�C�Lb:u����I�q�������������@'O�/{+�᮸S�Z��F��u
�b���g��� ��r�Yq�[Mr�J�{^��7�h���]���C̬��V+'�ׇ���I�����m=����n|�#*���C�x���"�ȆU�����
O�v%����4�����M����f��t`*v,"B�Z��NF�̮Q+���i
��fH��rǫo�p1E�[���k�$ΫoY���Q��o���Dh94kR�s�~���K ��G��x�t����J�(}G	�?v
r�^�d�/�lа��`+�$��Q�U��xm�y	$,�H| �yz;@;p����^xI��a�_��^s�_�D�{X��^�1+�[��0PO�>�ep0�;�S�I�e�o���^vj\�RŬno��_p+=��aT�7i���ҩPt8�9h���`�FW�R��,0�9���wn �é�����-Ŏ��P�1�v�[����C��)^����:z�'�_�dH�V��l����^�K*��S�z`�ṙ��8�PQ��	�A`��3{<�(����������v���l��>U�����>L>�sG�.�{�4�V�z��V�;M�
|�§͸��r��K�/��o���M�ד�U��N�����po�_�����4���.���?mR�-^�fױ(����Bk��u>��D,���?�
bY]��F,z�Q⢎��B��D�F���q1�ΣM��+�\h���B����"�ܣ��X�q���oL�.Iܨŗ��ŻS|�7�!�(�g� ��)�I5�ڦ�O��H�X���Zq�u�qA�Q���0Z�
& ��q_j�J뗇�~�AI�a����IY'�"�5a����n�Ϥ������b��~��tCwȞ2�:��S��S��_i�i���@�Jߍ���Y!h��N�7������Y��
���$u+���@�w~W���AT��6S/c���l�"X�Y������R�^�������q�}��&����Uw!:~3���R��B�O*m�'�_�I�Y�Ib�_�T��F����X��@:���O�L�� T~�s�Sw�q1��b��YT��"ԃ��r*�s�)��n�5Cq+V�,����N@I?F<9�lҹ�����t����aJe�D]������|2Uo)sYO�A ��������� F�y�I�I��^"��Ľf���m1 ���q��S�%EUOZGZ��F�;�jkpωP�%`I�M<�	hjy����#ǉş�@m�}���쨊��/��>{�.�/&�7�Ԛ;o�$��� ��,E�T��k~� O`x��J}�f%�����;z�Ol(�j�t�2�|I�} �d4)4մ4�;Q�
I�3��9}'n:aXex]g�d�mNT�qx�����;/eV*�Y��� S���+�C:<�V���.@��Й����������8���W1a���q����_}~��`��>|�6��׎U���FGY�1O��h�VwT݇��ȅ^�b��o�d#Z���0�휳E+�� q� i�C��}���p7/<��]{�+3�F�ȼrG���s'������&��jAH{�߶�G�\2����0�3R|(�b��TsJ��5�Es�c��ir���r�:/�m�y�J�mS�jJ�|c���F�ޚ�xV���;)vE�f�8J�*o_��پ�s�1�)�[͍�DK8��<�*�H<y���W�c����<+�	��a��� 3J��S�(v;��)��I�rL�&�����U�)DT;�%C�%�7��j�����%��9����r�P�e��b+�j�����}x~�șH�&�AK�MP�u�N3tk��R3Y�Y��~��=3.��?c�$Un����������~c�A�qw����F�h*���.]�������z�;���|�P�P������I>]1ӣ���t]J�$K����ᓑ�%*��f�-k�f��H�0-�':Wlf��]+!��u4����ڻ>5�ae�����F�<�͜L��1�o�,��.;��S�~��3�<僦����@����Ly��w*�����Q)2"d�y>��4apG4:
��O���F�� )q�0�̄a,�,��ͦ<�?�A󉟑Dp������oĸ�gLA�>Ȥ�Fl�X���{{J���^��afe��]�	j��l��E��>E����h�ڠ"S��u!���s�*��*��LZ4S��O���݃F�pp�:R��B�E�{�*L|�lQ�}:S��0�{ǂ1����$ XF���ђ$��`�e,ś�Q-�b�bn���S�cFDʼ��ĐE�	��x��wX7`|�����~������Y���Y���i?'����K*O�澕~8᢮��h_�I�h��8>y����e�a��q�.���%ts䅚�VִTb.����v�e�(PbL���^+���[��s4j~N���)����Uś�����x�F�������o'�������[��|%��N4c!������p�0.��ɳT5� �Tb���Ý�'^�A	!Oq����S���鏓V�
܀s���V��D8�P��-�}�����\Չ|�O	P7�g^�_}�a����,��w�E���i��"ˋ����/*�����$���L鄅���#��nm��b�yIb���L��E�������Spmƻ.����5�$��Rb��iA��c������
�Qtw��ʇ���RP��@q�	K_����K�յ�b��H�S솖�̀���N�=:�0D?�.���(V廜����ʁ�a'�j=�1\�j�$�@�l�Q�ݙغ9�lh���l�U�V-�����9���w����/�3���ܰ�!�O	i��a�HE��_��u�#�-E=�����D+���e|�Fw���R�,� C)͡|�X�ǹ��V�zʂ�`����D�퓦:�+hӬ1�����?��E��K͌�W��R�@1�R� �{k��ܼ� �KS-�����Ȥĉ��uZ��1�1�E�
$-�]����ϥ��V�	��1�V��{�JU\��ˑSM��9?�lsw:���6�Z�%�W���	���q�Po=L��ݼw������\']Wq��/��@�%��\�3F�l���$��pHQD���m#��Z;L�n���}/o�}؋�8�ˡ!I��l0�DSuv�\Ϯ�Q(��/���*:��]?B��|���	x|�ꉋ�)���-�|噍�f	�����T�E=�Y���;���3|�v����õ:�R�]7)��y�k�F���1�@K3{%��'2+�0�����~鏏�=�,�&�qkm�Xy���*�r��w$Y�3�������J��]�zFX��?i����a8�X7}yg��ϐ�%L[Yͧ��ˠ@L(1�]R8�}����P8֋��<�7K�����B=	���{��!�ԾD	�ɼǖ����LB2J2���ƻ��:�'�6�;�@-�ncw��♩D� Ӑsʪ��R�:�bCT�Rӛl^��X?��O�U�7�+�x��Y�Î����=S���:�'L���� e��=D�T����s�XT�c2]�]������@V۲͸`�o�U�&�eOy_�D��J"�	4�YaB/�ހ����0el���x�#@���԰�ЃfZv�LS�}�p�	���@ؗ���"t��� �;3Pu{�F#���;��1>���X��@P>N�"��ў�8��&�3�Ej�^�q/��v�پ�gED3�3c%��� p���7Z���o:��	M�m�单��p6ٗ�m������Ð\F�F�-U<e�	�L�{������1����M��;�II� s@����W�g�f��@����'6����qǹ-^}������(q�	�j�P}���̥M�� a�����[ݰ�6�i�ڢ�ƍ~��|�H�޻?�m����.x�Cѵ!og��;]�,
�]���My��Pd���#��Xz��/F��
/�֕��B����^�bcK���&����M�5�4ԩ�*T	��ʼ5no�R^��Z�.��|R��%<^�`>��]U�����P�8�e0J�٦s%��{�t�\��f��J��8��d$*Yu�8��I�%�����6���=X�o
��{�
H���*���)~"&������+z��61�&S(��N�k�b2�k�����
=�*����\̓�v��>�X�y��WrK�f����{��Qq� >��{m�⸆�(�_��ɪ��M�$�aDi£��7<�IZ/��;��\������IAc���L����0ӹ}H�]������|~�Q�M���n�s�y5��N�U�HV��yW�Y�#ݼ��FZ�Q�a�bGd�un���,���I;�X�����0C�&��O���<-E��V�$��
�j�"D�Z�X{,i3��7MS2����C'L����"��Jj�q��8���)*���e�BQ���+s`�/�X2��S*�s����d5nO�-j�Ck��f��$�lE�I��� ��b���S�zE1 _�:�V�����n��#�S6�"
��5)仴Hu�5�~�9���������X��9�+}!vXr,�n�!��N��!��en�����S�l��~��\W+b�?_q��+ܮB9z�X�k���W��I6�v����{��g��Չ���r6�wv���@aũ���8�>G��Ƴ�
��sGs�ѓɜ2�/��G_��E-�?]��4Q;©x	����1�7��80|�%ůg��tbk�?rp�\x={�3+.�Hf�b�4��Qv/{]&�MK�	��r cq(I�9�>��x�J�`!�+u�"�"&����
/�mKkZL42"e��e�,ģB����מ�v����Pߗr���+�~�е��I�w[g�����T3���L�	��<�o�����}gͳc&��R��Ϸw��Z-\���{	���Y�u26q\�^7bBg��E�O�V�)������p�΃����k{j��|�N*N/�+�%��ϓfח;��{m���D5p-�EB�L�j��.{��[�4�M�l܁meĀ}��"b����s�N_�/�_m����a*S�2K�q�/�����R��=�9$�l>9�P]K |-�+S��U4.�1�g�,��-df�]>&�%�{>�W��&Q}@1Y�"�p�S��S��/50P�q�j)�ٍq�w��p��ǚ�#��%�s½��.gҫ-�u�T2ř�窩�,h��ؗ�v�����d��+��}-B	��_-����d䌉��l����\�2�GD��_���Zo7LF�*U+��%3����@�Q~I�(�֤2,����[�����=�U�+k�֗��!Ƅ��"W���"��w�a���5����ӫ�>�b�x���E���>���@J�%���U��	S$��s����:^P']#�<e+�H(��3��Si��DE�Gdo%�����2"i�U3+���.b*��K�bˈ��x[�$�!��U�a�9�����O�V�A����@Zr�Y_���zY}�� pp*Qqm�5WdEO��j�H,�{���+�����u��&Vr��v��倭6j
����$=�,��P�s�7 <�Ѱ[ھStc������Ƀ2"J��9b9d�� 
��%�х�
S���۞Vآk�r�r�������0bt|ȗ?rZi#�_����!�7rW�LZ��ap0���#��=�h���qS&8�r���ۈ^��gOr�	=�g� ��٘�,mƚ�Ke����0g��b���V�4B'xl�-:�Ob%f>�C�+]ƅ��R�ˀ���~��i����v����.13��s��i
�����u�{�Օ��_F;F��4�5Ƚ�&YV�ѻ̕oґ��ں�ѯl�+���'�]�o8��`����f�M��$�٪q�o���C_k��-�o���u�W��R��\*߻�%��!����網�*�!w�]W�	��|(Q$�k��Ŋ��w���e��ŕ�	2đrAz�$.!8>�yN��q��>���]L�:�u^�������:Ԧj\A&�9ьɠu�
�-׮U�{�UG�*ꃶ�D�ĩ��Bެ9��<�2q7�qm�V~���m"�΅q竔	#���H�[z���'�?�
�~�����Vp���8��+�N����T� _v�4J7��qJ�"m�#�B�u�)Ĩ����]�>�^tL>H]I�m�Z�C��ί3��|H�@� ������LZiy4x�l���h�/`UV���.��>�%�ƗY��2�oܬN�o�(\������p���8׽.'�b85S7		�0�L(Fq;&�Ti���C�X��Lj�\�G|��
@�������$��&��������!W��W�q���CD������!���S؄�� �!oM�0��_�qBԑ*�0��+��q��7w���+I0Y���.#��|�KW>O(4���*��l��$`F
?~YP����X���4�t|�@Y&��h���3g��������[d]�ۄ��-�wsZ!�9����<�鬚�,�$�ۭ���8�O��l4ix%f�E�ۢ\0��p�p���
�H�ĺ��n6��D�W7E!�PBJ�����{Teg���K*_=��?t���5�<g_�L&r=m���=���r�On����͗S) iPW%3�#!���/� �z8�}��T�Hu
-��4<��?���o�$�O��U�2j:�)�Y���f�>��*p�)y�HPݮ���oF�|�n���es`�8�ʡw��sWy��a�؎�� �q�ƹ�`��
5D+F�Y6r�N7ui������ʛrxCx����u6u�`�Ii��z7�F?&s�7��Ӹ�n��`@;C��D+'/���K�'z�+5�����@�R�S!2+���v� "egD�ՀC�{No��^�y�	�Idf�hU^��z��S�H�8,1M�%ͯVbO^i�%C�O���2���|]Zo�r�ϱ��R^����M��3%�7p���JƎ�:P����mO����v`P���	���9F/=%�_n��~�䪡͊�1/-V�I����Z����gw��	���˔��P�s[y�S2zç�*�����X�j��9��ӌ�jI��(g^f��>�/�|1ė�{�����7����O����T�d=�=�w��ã+�]$lZ���2����2��g_�BȉE3���{wt!D����d��������.l�!^�s��u�9�b4z�kmZv� �w�- ��6>��;<�`�VDX�|ΌX��|AoJ}V��T�X��ۧ����)��C4��!�;�C���h��j=�44<LU$>�8�O�ܛkBC�|oy,�s_�G״������K��!��]�8,��	 ������]ߒ�y��W5S;Us�̱���9ݽL*F8u
R�c�.H.�h���Y`��=2"���W�,hh�������Z ��BM�-�q���ԡ��<�������ۋ�ݬ`R�o�`���7X�4ނ*�S�`��R;cQ�mB���H��h�{-y�y� 3����jB�]07�)60����%m/BхСTc�ԛ��6�:$�g�|[�Bn�R耠H���:��88�?��i�!�c�ޞ�B�?Z��Ю�A��6X�nˡ,��6�_����&q��󰊂���!��}yC�=F��.-i�#˩��|4G�����0��yRi�?t&妇��:x%O��q&t�i���u�I��i��*T�4��z.7K.�	����Va"�lj�Aɢ0���� bH�Z��h��f5~of~��8�@C���!�N�J�n��Ӻ�w�.~�v��5/���.:�Ա1�Z�+ڠ�?`S�� �v�Cݗ��E:��,�mt-m�R�y"K*���������l�'42����![���T��*�.&�Z����J����������w��b�?���m/m��q��@Y��+��n���'��e'��<��nW�K�Xc�CK��S��}B���.[>�q��gFk�W��#�!#1�ٚC��q�>�;ҽ�Y�ج�E�����2k.>=H��2
vb��*�>7�%��2�	��2@o��fG��7�//%�yGW
r�jW���~T��Jnxoxd0�A�(_�,���ݧ�j����z�ؾEA������h�][��w4 ��}�,��mM���no����ͺ�� ���ď���c�cK�L�w;�ʆ�A�՟���vSʄ8�Z��s��w�]��>.>;b��U��v��n`��-�zac/QJ�|�1��E>Ԗeu��%���=�."Jun=,U���[B��U繺�έ}\��_�l��n�d�u�(�8�5aپ^�ͤ�W8�e�Ü5�G����$'R��Ow��u>��ñ�z��ng��k�g��<�T���}HWpu�wJ$���:q��tBe�]v�9W� У�}-l���Gcُ ��H�������[���9�X亝�����u��V�Zy�
��	P�^�l��RB:�BuF�� ᕆ�H����~����ʞ��p�-Q��M��'H�)���d.�s~���?�R`���>���Q�@o��x�`E}P�.�iu�ab�+&3������݄z㢪��qX�F��!��Q��;��4�O��Tߙ�M���=r�O��)l���~� �.s/�?��ݓ��G���r��x�7��`�شc�_�M�i%�d˄i��:\2s�� $��sڎη����B�����<��I�����W�/����v��6����.1�:'N�1�Vڷ!�o�b��͆5���� a<E��S0[�&x~P5V��Q��غ�zO�zN�TE�qcVݯca���f�Zb�(�)�a��&�]���V1lVg)�W����V����aVcT�5U�ֺ��6�E�F�F���2E�HJ��IWx
3aT���ڞ�fvQS����3/����u<kH�x,��e׮�x�T$��Fu�j��Q�lȘoW��R�%�s��`�VyH�>%M���I�WD`ty��]E k*G��%q׼e��T���Shw����av�8�>h۽R=��^��H�~�2�B�b��a˽�?ˍ?k����@�O��\�m"�p�oz����=)4(L}���[�5�gmm�h�Ehr���l��> �M�s�����h���d��!����I�P���f�B4)g_s�����H7!��E]�b�O8<?3xM��]_<3���	#����h�,Nk6]5'0�MzU�����/'����},�˧��O�D1Vw��͵�G��8��)#�Ѳ; �5�� ���^�'����"��%�o~&��լ��yyEmA#e*�1��h����|�B�{`eM�J*Y/F���tis~*_
�J�~�l&���=��Q̂��
�[����Q�u�(cL�{'���$�wġ���n�.� �2�pZ	��Y�P�r����N����-�*�\��d�/q��om(��F��J��/�Nz�=�-YtT4��?L�`&Ҙ1Z�o�N�n��:dr�������2�)���5�&f�N�2�� �*e`c)���AY'����A��Nt�R-�_{	i����X6_��G����,`�3�[�c?��SF�}�Sà@���&���PF"g����޳�ͺc# V�ި.�?m���8�ڦFed8>'H�]�]^��D%ㄏ.��բ�rK�|�`�g��e��9r��ӑ��2��C.��XS���Bb)�f&����8L$4�$B��O��S������s$6��N+%k
m�+/����:Ӱ�*- Ã�x�q�pZ�4q*��;�M���ۭlTCL��D'�r�7�9<3�}O�C���ዖ�9O��:]�k	�Vj���m��� &'��wsW�"���Z��R�.����]����ިU7_S��l5��7Z�'ⓛ�!���}���C��?�Iz��?v �#l���beܐ��p���)hoO!�l��7л��E2c��w��=عe�
���=�C�`�s��dl��=�ҷ0Pt�^b��>�"f|u�69�Ÿ}�(l���?��K������HN��;��[�׊�Q����yB}���ˍ/�;t+��4��|L6o%���,���S\��v�!��I���Ēb.ø!��*�O�ڹ�E5���-.[ٌ��ܼ���蜮?�]�>�5�(��EY��X�l%���x|6�X�c���|���T&�0M}@����7��6�R.���6u$UZ��d�7Ok!�w��2��5��E�##m�Z� ���FkK y�]O7���E�Ո�@�B��:�]tR�@]�6�"҃C���$����`-��yj�ɿm����~ݛ��������hi�a�2�T_�^��Y�������䯂t�顷AA5I[�mb����� ����� �	~��'z�X-̺�n���N-)ٚ/�A�s�������?��q6tp����($t�ǲ��&���eN!P�6�M���xO@�8�$qd�����`h�o
LڜϮD��3+�b�����w;�f���3���ċdݢ��R?��K>�&nG���b�*l��Yi���Zj�龾p8�����7��I|�����*��J)/�B�F_��{��2M��v}�H�@�
�iir�<��h�<��AT�K�x�-g:z���Rtx"�5��
~>�vnco_�5&����xDs/��$h���F\�΅y������5!�6X6�>5�(
�/����u��҉	E���~�rB>"!���E9����G+L�f�KDII�Ҝ�g��q�o0��*?u=翆�H��[��V?�I��s��u���?Rq��&�J)��H���T�-�8.eo]t7���9|sbb�L)�����'�N|�e�M����؎����K��D�a��<m�L|�)瘈!�+_U=�@�QѴ�"P��q�;u-{�_�u���m��h�[��eR������U��a��L�u�p�/3I��3le��RFZ��rR�4q7�c?���w�8T�˵L�~�@�������5l>�&]��|U�-k�ou�On]%Dm�c#�^�u�>�4��i�p�����Z�#�]���$_`h�J�ց�_�q|a���������p�<�<H��eC]��xdW.�3G9�èŌK��8eO��>i%�+��q��Ѳ*��8��9��%���`���{Qݙ��f\�T����1^���>m��h=�J����b�y ��s3�į���>���αw�q�d�)��-|�A�d�e=s���SZb������Mt_�H� 1j�{�����յ�Н�Я`qMD�}+����d�d�^1�@����������|�q�u����V�S䨼�;��&�,��?~4Q��_g�q@y&zb�L�Y�<���g���#GuE��������i�	�*S�����٨)(�wz��'nB'w]�n��$��5��	�0��‍0��O�����1s�?-P�>�.E��E�XqNL�=�'/㍵�qW�qt���Q����a�������$�3�4�ټu)����b%l�K�+V޾�&�g�6n]ַ�ӳ�1��U�����qE���?���������@��(����u����2�'cvZ9�/�R7���*�f���"JI�����#>];�/�>�o���^q�)D�J����mO��/K?�^�i��4"���d����u�Ҡ���--�NE����[Y�,��{a5��V?�p��]�eV�������M=�o�L0����+~�O�z�5Y���\��"�������ֶ���3_�g��qi<���gC�v�s�$�qM���3�T���R)��J&��w	�G�`�7����R<��N��ݤ#;ɪ�&��j<lB���Ƚ�	H��y��|"�t�qh8NHA}#ϙ�Z/Q5�{6Y��Aިǫ7Y�l�H��:��d����K
I� s}+w�4#���"��c�*>>�G��}n��`���"��A��B:���PO�H��)��M0� cQm��X�v���5�N���Ȝ��H!k�2�vr�A��ϊ�?�\~�ow���W�pD:�}��p���u=ꍇ�h���TAA�$��P}oR�յ���^�,�����
`��������s�Ը����ټ��!M�}q�����[xAG�Z���s �V�/�˗�?{�}s�'fOSTm�%���jeJ���
p����	N,�����ʛSaХӉ�@D���(���SE�{�R�˹��7cb;�`.�_��Eڕ��B�����ҽV�{���Zw-��;��Ƶ�F�v�ݟ&|��֕��(T�J(�&,B�d2�H���eJ���6PR��1���^���H��Mt9R馀�G�WqұS����yr�Y�@�x�c�G�<�+� �P\T���7G����B��<qC��}�~ۍ-$����_;�\��Y��>�J!�B��h�ge��Tj��o����+ϒ���K���sOA�M��b�߇� �i��x�
�	����X��
3NA��XC�"�ˊl�z��W>�@����J�R�`��㟁��z��T<ҷ@��v�bM#�s�	^q�FA�ߘ?x����6���ո�͢�1<�d���|���'z�ۤ++�����~������� (�+�r�~�T:�X�tc�R��ݫ`M�]�ao�-ɵ�)�&jO�W`�֞�!0��v�(��kWCJ���M�����W��f�Y�uw�R�5��нs�^�Q�{�X^-y��1c$�?�ר�E�a!$0��q�Y���A=.�����G2*��5���ټr�D{|=h��v"�&��_g{��׏x��jF`��>c��8�ς�d�{���_oC���u�U���s�`!^Ǣ�b�������r�P�컑�߶�&cG綥hyT�m`\+�_����kj����Gb�䭭=RAj�h�?u���	������s�:Y��\J9�n�L��q2����Ao����_��}�����Z�)�iU���` a�����_�S��k�^ƪ�Jf>��6yN=��5l�@{w���Bli���3�q$Ė�	壡��k��x�����e~�~�Wji.r��`��f5V��O�� OO��Fw�~�P��'6T�5`C���x������~�*0va�౛bjL`) rXJ�T�ᬬ�=X��0Y��R��b��B�c�h8�35���w~H���<"���2,�����LQs��W/s����� Q��¼�"�y	Jh'�:�}F@���)�}ʫ���Z���-X5�vm	+��"k��eVO��w`�'M���栁����|�X{�o�t�0g*ѵ�����/ �M�V��@�T3ʱ"W�N/d`N}��)S�K�{��E����e
����Xg,P'e�#���u��K�$�,뫤�?�����D�Z���|�|D+�,K׻F�%�Q�.+C�8��	�#�+8݈�v�P2x��~t��"�đ,릣:E2���)H�1�"`#Ĺ�U�u!��}��=�,;B��H���?͘�Ș�x�D@޹��k��G�c�۸V_��d��`p>��sX�����eLK/�kˑ1;�Lۯn��:g^-�����ﱦ8��F�4���\ �����?w�D6�w_\�1�pk��K~��'��t_��\&X�n�:	�x�b5�b�~�Fx�V6a҉���������d�� ?�FvU��x+d���H�f���&�_g��/v
���TkX��[F�z��!iu�}�*f"���6��{~���ȓQƧ4���a|!�o�E]2U�+.����+W�|��/�٥�yi�1�>��ނ�$�?�ῄY�G� �Gb�����6G%\�ޔ�k�OX�[�m}��p{�+I�����"�^'$;xl��%a�h�#0�X�I|�/��]�G��A١��(Q���-eEBm8�-��|o����2@��|�.�ɠ������T,h�18#��\�9Az�x�N�4�Ě�[�;2����}b<x� /��^���i�M�>��2�ȶ����6�)�e���ɯΝ=N��%��{���Z���NT�d��6������@�z�E'Wo�ъ�A��3�y�a��	�E�Of�Ѐ��� �����Ȅ�ٸ�P��^Gb�$��Yj�W�ҷ؅j����k��U��د�g��3C��G�A(�~9�^��Z�6����I���o�)>[��3�gr4c�@��je[�;�©���?�ى���p��IR3z�-{���R}�ۻ��م���vfMg�z��ގyP�os޺��o����?i�F��|v� �E�@w=y���zR1�S��t�J�6�0=%]`�N�;a�0J�c�+�����=)�?őw�I�>���0����$���Y����r�-�i(��{^mla��я��o^n>����&�U�`��h��ݶl��*݇lj%�(f�����#B�ѡ�d 澿}���S���6k�r��=�v�L�	 <+�M���J�m�:��FO�u-�II�߿��voc��MY�O����cIN1�t��0���I�\@gό;��O����c
�����1�D�J�Z�
�H1���_[��W8w\)&|ϳV������}<���.LP����=�Czc�`L]ب���%U��r���~Z� ��qC�]	Ɏ�>8⻞�[�"���-���F��x���	B'���e�am>1r:���k#���?�'�q��o(��q��w��^O��$��~Π�Y�72�d� ��`�=��U��γ!�N�E�N�F9�����"p�޼�(�C������e�؂Di�l>�xi�A� �.w~�z�`bG��OD���r��{�`x]��{�4Q@�sJ���΂���Xq,T���1�FĬf�o$�Ԩ�>FI�o�n���Ƈ�.�τ]�����ƌ&��]�E�iu�c)�ij�N�oJ.*$�EK��ju��e|�ؒ{��'��~��������co�p7�A�XA���������Ĵ��s�G+�/mth��g�w
>���I��>��)��J��wbqb9�")1�K�R����2>`��H �l&�h�u�(��R�B�P�4��@/�Z���AS1۝�?LPU���*4�b��wQ��y{C.�oc�-��dH<[�rP��hF���F?��	X�9*��>�RP:f�e�z�T�Mn�����#ҥ������T��f��}���oAt��qף�@bb_��$Օ�	Ĳz�u�&`ėח��7�D6��!�����W���oo����_=�ll]�F��m��ӆx8��^�����v�UQ�� ���I�_���	��U,���K)¿��m��2��5��y��@ܽZ��F�:"��s
%n�NQ]���\��2�X� X����ý��n�K��f4щƿ�f��U�����Ņ�iLN3��i����ڏl�r���	�h�[x^cH��JL��^�h�����t�d2�nJ!��TwK*t�7�����9Z!�P(�Zǲ˦A���3�W��s�i
w��5�N�ǟg�� c�Q5ǂj���KmgΓ�_~��9�����#m�[�%� ���G`b�u�����/XҜsޮ��b��+�xB&��B��J��C�2kٲG/G�&���q�4�`q^\d80�wA� 7�0Wۉm��N�g��oA&v��?[a=~:���Y���L?hY�T�V�'Ö�T��W�"�۲J�@J�IRd-��u�Z������$�PIT(����HV,A �ܩ�Q)�2�!�J#��Tڟ`��Quxh �(��LO�s)݋�?�OA>��۴�K��0��b�T�Ϲ"hM�(�q����O��pXC��A@�3�y�/���_�{���S��I�ZA�O
����"@z@��SS;��&G���'�U��*z"y�_V�X��ڌ+��T���k%9ϓ)8(4��S	��5&�� �N2��?��?0�8K��g}��,��HM�M���P<�쮵�zG����vG������64�!�.ۓyr�r���Z�W�P��?����7�Q`�/p����%��S��+���+�?��$��#|�򯰜$��������t��V�i�е�$_=X�^���S�D�L��H׎K��Տ����;b;���^� ��>�_��~z���!2�̝���G/�y��:|� �Gw[��<�M��h�4��Y����,c_���YȮ+�ꌢ����L�l 믬'�����Nr
�֍��k4?/���P�dhw?uj}Y��M��"�_�r?Ee.N��L�=?T�^��v�r#��8��=�=~$�a��S61�et�$O��_r���y]�ڀy��o����ﰩS�/|��Ĩ��Z]v���}-=�a�t
�5ձ���ԵxY�vl��.�_�����[4�V0f��v�8��֟����/'#�~L���Tf�G�{�ec�!P8�Q�����Y���B��O��,pE�����"�N壊6��65�$6{�~�2�l���c>�4^��(¢�_��+����ާ!\�d(�u�Yʃ��Ť�r%&P���� �zȰ?��َ\�uϴ﷝�� EsJlQ˷���/o��5'����P��6=��2ZrT��>�8Y��x� Ɠ_��e&�'�/2����,d����̝d`5����a��n)�ї��-��،g��P���k.+(P���?5qn�~�dc�N�].Gc�c����T�L�������%�\��
�T6m����arC9��\:P��.z{��s�tp �����	
u�ϵ����d8�� ?�K��b����9�w�]
�
�8��'7�a��C(L��8��,�u����f �T�9m�]?;d�F�&�4'��cf�_$)N��-��d���l#jat~�j.�JןM\�~�����/��1�� ��b3�8�T$a|)s��:쇅�DD�Xb���?���L4sAh�*?�����>Pm&\�����ϐf:VM�G��22T��rը@�M A*պҝԕ�6;�'��+��T Z2���-Ѓ_�Z���������K�M+�Q����C!Z�؝���Č�Y?�����h�Uk:����S�`T��G��yl�4^�X�?޻v��7�F���i�����${�K�,�m��,�#t�����s% ���W���C�O���HJ��B���q�����$�~�,g�,a8���-P'��F���Fd�W"��4+�r��/��%���� ����BWh
w#�BJ ���􂣭�͟��:��.�X�#��>-���?�=w���)\�͒x~tڂ1�'&�䖠2��U]bհ���c�+�M�q� N`�:WVRϪ��w����8N��2nd`R�E�,Y;�e^�&%F	5{��'S�J(���S~E�-K�c3w��I�g]*`���"�o֧��kO���5:�$#����	�a�"׏"����ͦ�O�� �Y4(�oPi,�W��.A������-S�k���g,)G 1_x��~3���� `���7��a5�����F��,�	�ˤn-�j�TO�
_�S=�G��$��N�F�A{�h�<��<��<q��F����\(o���ܸ�d��&W��uE���?V(T4 �vJ�=�?�=���@�&���|9��5J8*-2#m4���e���9��r�6���C`@g�OG-t'K��l��E����]0� ��4M�c�W���y�J08�2s#<�3|@���8�>�vF[�0׽[uh�NX�p��_�I�d�U@���W8��x���d�#��Y�S�p��-NQkh|)�U�MJ�J�RR��k `��"�^����㲲8B����JB���BL��m�X��o�B�!�ϑz����1�!M������͗%���Xur���-�:��J��|�]�u�T��b8}��}Z�7��߲��Ĵya��T��_�̘8��ӎLÅ�!�S��*�?���}ǳV�Q���~�P��K:W�b���o������j�ځ[Mq��-ݝ��8��S���+�U{g�Qr��v���r�N��zsw�[��yid�\�.�X��S�L;��'˘LQY���{r� ������,�LJ�	x3�0]R%iX ږ��Y]�%λ�8{̍��)�E��*�����Ч���+�K�m
DZ�-D��䬅w���|ӎ��8�b�0.�,�~1Ȥ.%e�A]��e���
��%�Ai7�g$XU��s+��~�( 9Ѹ�嵔;��� �Jm��j��J�MH��*ч��%^s�F	��8
���Gen�܍�l#I-JHy�Ⱦo'�J�'<���h�����rNj,-��{��A�do��L=��bT�?�Y��FO0��������~͐�<a9����6��oTPǚ�%�V�h0	p�� �
�1ʉ��ƶ�x"o`C�|��Zs�'6W���D~�ެo�NfD��X���_�0�w�ظ��V���{U8i
�ٗ��idn��xG�2{_��,��A�:c�Rx"wo5S�E��k&��.]�����f:,WG���4�A����)�꽣и,ݐ� ���G���(u������������F�����I�!E��{3=T�>���X�9K�b-w��Z��b?L�)�׀�KI��>Hkph�7��DSl��u1��nv�z�����$�;E8��f0㚌	၈VB��z�0	0^�RZ�_>B&���5y8M���Àl���&$F �� ��}1�Dx�&�Y�P~��P�L�#Q�������;�}�4��>�;�~���&Mwe�ܐ�ˏ52��U�D�@�;�u�'F_U��Xq샗Bt�3X;�Yݖ`:� 0��~��	��0�q`�V�����BŚ�3�+�F��H*L[_Pu�}?79�~��lo�xL+�q}�L�P7��A���\����sl���T��jv�����V��C��{���|O��*�y|f�V�������\6�z��j�1q�V����K��x�˚� �frQ��.7|�éoP��Nv�^��o:/	Rp'��w���".�DV��J�5r����/,��(ܢ'� �ۍ�ּ�0�Y�߄y��#uR`#g���G�~W����p�e��Â����J�GM/��A�P��^�l%Y@����i3/L��ݼ7�R����z����<R,}]3��K1xF1\I��Be�~�+͔��j@=+�Ϳ:���g��-��c>�t��~]U]�؄��9���/���vt�_��M���i.D͊d����T��7ܖ����<����
W�����s��As2Y ��vOQ=��m�>�)u�����u���+�mw�:0��sR�����n���V.�A��r&P����4�8Ws��o��3s�Q5�n�@X�:J�ac^������~�@� �j��`Y��'���__4ʠ6�[]���z-%wD��1XI����|}�HҬ �,�=\|Ǽ|����J-���,	��B�����_�@U���3�'"�$�,F�`�)7��1Q����$�����������}�"β�E�V�@�u��-Yф��q�mk $5$�1�H2���}Ԥ�I�$x�pq�2Bt/J�^�j\����S Xj�M��g$�G
U4@�S� �>��%�������g����� ���T[�lD�j��Su��~���P���Pq����9=�uIFqj"��mk��T׌;�1��	ٞ:�f��Z ;����B�a/V#���yZИ�=��\3���3�5�J�)H��^Y)��wLg~�T���(>||G�hʼ!l�H�d��1<����G�����~���X\1h��	�FV��CiF���dD�ђ�D7��(�H�����X����E��CY�ċ�QMi�0��:���	C�|.��ap��vj��t~���Ph�l"�.k�E|��4�k����_�`�� մ�wd�Eg�#r�e���d��<��dֵ�����ǲ@�jP������x���^�QF4��*��k"��~Mh֏j,˴e����
�-��?u.c .r$�Y���_IL3l2��r?����-��
�u`c8¤,� trW�\6�²�]R�\hf4;�"�.�1�����*����s���ІM���\�@��{N?��	�n�~����������������}(M��rj�h���[US[U�H��I�b�(h�mM�WN�	��ɜPC��94}g"}�Q��#v�ߟ�
�����8ߍh�}E1@��(��J�'
W��t(����v��R��<^ûG*���2�n��{�6�g&Nr���A
�D<��?��^xBp#� �Ҝ�a`�����2DTl������������j5��xq�ؼ�̷-�|d#�'�W���pw7�Q��j]8��y�HxR����o��վ�,���QUSN�0l3Q��']�ٴ�S��O����^5�W���t:7�fĨw<i��<4I�d��S�������"�bp)X�S
9a-m�C:�l��r@|�F��㫑�c���i:ib~r���n����3Y��&�Cʓ�-��7P�x�2o��31�U����\-��m`���'���	�:��#u�
��q	ń����$T�ЇN�~7b+���������V�f��CD����(��Nk;�U�KQº �����4�9�&�M��M#���_�i�����Y��qƳ�`*�w~ ��`�aBU
��=Mqk�A��`E���oM�J��GKO�fFj�&wb+Պ	Y
T&�Ƈ�=�D��[)�	7ad/��R�7�����i�m3����쳽P��R#���tC�@v��w�	�^�TX�V�H6�OV>G���͋�@7�5�U��EZOխ{��Y�Hek���0:{�p��&�_^ �鐸���>��$&KjG|X-��@�>h�[�����M x\0S���1X���vV��� �V'�����6�![�h$ ������V��r�/���~`�G�p{{^2��Y�:!Kr}��	��5�7J�e1�q��>����`��|좡8��jp�QQ^^���#��?� �����_��;�ԙ?��.T�2����B�$����\�}������q��FT<w�ɎU>f���%�f�)m�i9��vk3��eti�FE0šLbY��o��*#,�t�`K�����w�E�(�0>����9}W\����� ��P�"C��c\f�'Q�v�������BBWC:�6�>�{��͠�Þ�Wj1�G�q�鮓ݯC+�im� �Q �ZD��:���u~��عA_��$���myg]`l꧑`	F��VAz�����5���M1��9r�F�貃��.Ã9YB�IT
�]�:�?Yk��):=x�[�$k�@�-������0�z�e$U��mz�uFOZ.����L��цH�c�ľ�!����DxB�2��[1��`��>'�[�h�Ǚ�ȗ`���3�~��Z��W��6������̘��H�H����:�8-M�j/H���]��;n3�!�q?�>�Z͋���������MP/P�p�񬿧J8���G��X�q�����@�Ӌ���g{�Ȁ�.4}�X�5'#�{'�c�F����t=Ʈ�Vŕ��9�<h�?���IZ4S�ƀ�]�g��m9�&���9d|��R�+�Q�������WG1�41s�[o���j�*z��WD��
Ǹ!�	�<�������Г10@��Ƣ ��8��Zl���X�O#�V2����ψ�)f�h�2X����q,��ѱ���B����hWR�i�9��]������3��ױ$9(Չ)Zl�E���p���p���0a��&��S��o��!&���H��#=�6d�ypc-;F�W����I�I|+E�K��I�m-J|0|rW8��7'*S�>i�J9?��/o��B5�U�z����1��+tq��|M�T}{��b�"�*|^8�:���c�����O�JE�U܀�0�t}.�K�#�,��Ä��v�z���e�-^'z[��b+���N3�X��l�>;�EKK�GV�'�|Vq����(��َW��:�P��v$��,ҫ��mz�|�:U�4ZY6d��̫�d��G���2F&x폧����"��{������=l���vVoWO�Di�ÿU.�g�/�Jaȴ9s�4�!� ��y���A�zYy�0RRl��X�p9�|_h�J��E�&�ǧ��eRu��EK�TT�t<�=��(:j�Dq'N�#`�< ����4�n�j�R��E'Y��^�
:�y��{�����$&'p�+��O��X:���H�a�\3�;x�w�,|1��\��Hr��qA��������v��*��e�$j4ï���}���b�>����^n�"�����F�<t=����шQ��������.���=]���`��=�PP��W��(Ğ�]r���en��Q l���̵�����3G����w��Rq9�K�����}�UAxg?���a?�U!��k��<�A�S�?*� /-�:k�G�� 8&"&K���۾�˞;���"�/;��m�!��?tT2��y���*��`I��߅6@C�v��X�ڭ]�Ş�|�,��L�Ҿ����m]'ŝ�B�ͧ)����5~�|��{�1�{��!���u��ʽ�jr�U[�����l�,rE�v���r��gѨ���	�vkcW���~T�fz�hN-�m�7�Q)*0q�w'�`Q(���\3@�J�-[�僽lNM��4b�ߍ�#W��vf �1��q����G��uO\V ��5u�����6v�ǰ�W��l���W�t@��24m���-cS+qh��kܾ��ŋ�����	L�^�~B�.�b �5)�帑�>�>,���MK��C��|#��,V�A@%~Q/�3�׃A�\A-Y�?Z��R�,f�{��@��0>Y*�w�CŅ���1�T���U��������F0Ta��q��ʍ�o�����	�9R<���6��?��܄Gh4���0p+��������o?Y�A�T!�\�S�z�;ÕW*<�1l�����������Y��GS���~�<o�Q�0�R�f`/I~#����_�A�9�S=ROޯ��}s'ǱZ�ة��9Q�=�]i����O�E~��QK�i�W�-]��D�9Q���Ev��K .C�J����Z5�
C�%��x�(�����@����+g������ֿ�C�bB�z�+�a͟��18Ioa�a�{b�OJ��/_��)�p��x���q_���)�D���H�*�Fģ(��n��:��=H���u� �;�T����Mk�^&n��������	]���ع)�e���[�_;G��1W� +5�Q3}ڗ�r����XK��c�?DT���i���7nUoi�I�R�2���q�%	J�J�|��Tߐ�C�it�>V��dB�8�έ��y������S�L �.o2&^�(OG�v�(��eM��~�87ݿ�������5�i��2��n�g͑ ���;�ҁP��e��R��x����`�P�0�6Lt�-�Lt$�M���*,���ݦ�.�f9��\cƥ�{}]�ߜ�w:�u���Uڙ�R�8YY��M��v&:n�]���M�&��4��?p�Q��D�?��x�>�#}}Xo�mAN�1�#X��/j2�F�,�ʃO\��t��TJUe�u	���q���Pj��UOG�%�&�#?�*�]J�cWM/;e��.@�Á�gM����Y�N`95��	Wy�ܔ�:��	Y��&u�1y߃{J�'�2�O;4c��U�Ų�)p��B��驅���#��-�E��L3�M�{nñxQzz��˕��_����[`R`�� &U=1��S{�R�fc�9b_Ioo3�H�\�־��u�o��8��Jk&�;��L�-{R���<�[%;���?��9<���zc�q6j��6��m�vۘ��ƶm�jؠy7�������d��[�>g��Y��D���&R^��W� �B?R+l�Ð�w�u�a��Uֆ�X��f1���j�T� l�l���	��ʉ��4i��c�E��l+�)@�]V��r�.�.��3������:ibDtm*2ڷW�:�}��Q���lQe��Wy���˽��x�ώ���_4Q�(n�3���:���]�	W�|m_8v����"�I�>�;N�e� �V=��O}�=3X!���F�P�@MO;�@?�l���:�5y�Q%�ڏW���Oi�S�ZO��ɦ��R�ߨB y���j_+8�*�juLrj�5[�zԆ�퉵S0mޤ�Tj�C�vQ�\��������;�FŌlv��W��+%��t��_�������������W4�t8�-�L��P�!� X@�r {�2ב���v������yĘ����o���!]Z��~vD���F,��FN÷�$|��-�>$RZ�~��H�w�4fb��OD6'�Z�Zj?��@`�jk|��������8��f�{zNd�2�������E��{�ȁ_���Zč����~ =��/;uz��1�Ķ�9=V�I9���29Q�)7�J���7��2������ܨ�/��,�'�-��$k5 )4���?[h�=sk�yK��S��B?-��+R��wi��%��;��x���.��\�7,��Z*'ޟ�*o��,�1�2x� �W�4�:Hws_K�$��;����L��	��yK��v�S���չ���I��HZ�(�i��Ռ���W¾�_h/�#x���D��T�}�ǽs����苼~�>j���P�)���A�v��r���y�Jj�&5v<�0[ۍ����p�_����W�-m��9t���5>ˣ�"��X�;B������wE��w}ǽ�mŶv�8�4���f�6h�-��T����Z'�qJ7�,�s%3�S-@�wP��~~]�^�&e}�2<8X�;��	{AP	����/��=����Z�j�f����Oz�M���~s$@�~KA�Eψ�ɯ��`7��7�Y ��N�j����� 3���T����ᖻ�"|�x�DR�
�hr>��tG�DI�8d���	!u���+��Ȱ�8�U½)8A,}�W�Y����;h��5���aP�� ������+pYS���c��
���Mg]?��o<�����-�3���������T�V��k�+e��Ӎ�J���_�������ޔ�@)6�'ً����j��� 	�ɫ ����CN	��+�R$�.��7�{��������}F�׺����7�����u�����C�fZ��3*��Ʒ��*wO�Dw��v��
��� �8���i���J���]�{~ m��y�,���� �`2�O3`c�
�vsO���&�b^�=VmG��'��QǹߢQnS[Z��,��!M	��n;i��C�k��i_m�myG� J%K���w;��K7X��3я"���Z|�_(�x�M����3����uZ�v]�%��@�J�T"����,�!�,+����K���u/-*���t*��a%ޟ�J�[�v*r�G:/]bk��i���O�6zLiM�V�����t�4�mG!���Ԕ������_3-T'==;�Ϡ��%"��R��Ǹ��V�P��!��>�u�FS��bi�������}�k�y����u�z��yv�y�F��+j5tn[�2��Ea�n�,������3<N:Z�O8�\��z��_��KL��9/C8�/OCt�|H���t�)0k�e��r
\��_��?Ԗ؟���*�,�A�nz���y��� £�ص8��{Z\�����-�(���ӿ����d�Z���7����j��f,^`ÇL�u�2g!"����n��� v�^g�)cN�R3�V��C�/G��>!�A��A�z��+��1���ȿ��,a��CEC�^po����3�~��c�+�[�.�������͐H�u�ߘ~��X�#�
��Q�� ꭭����%D廧�r�7mSg����J�����A�t4���˂����^��Q�J����ӓ����;���fBٛ~��I֛��"�E=6X��~������m���;�Nk:�bt�[!{눛�T�R�����`9�h���,B�̻��|ғ]��;�/+���=R�cI�x�o� ����a+f%t@�;U���/�S�WTo�L����(����ٹ���N���[9˯�}������R!�?ɩ7�����-��{/�z\�/K�|��X��}	��eT���{搑�P������E�9u��]w�r7,C�Eqn�PLj���Gh�����x���Q��BxUVZ?�3���_\�ϭ!rT��'!���ż�������rY��у+��7��iyx�T3#�ӗ�o	��󰍜،�H��J�p2�W�/���P�x���ޏ(/M ��O��R���z9�� u�~���u�>������AK-p)n��-����t����6��sj������.:���*<�r�B���@V3�����4<���㺪����ʒ��m�H����O�	��u�� j?�J�|Y����`�l{{,��	<�U�!�&���RWKI�;���<�6����x�ʹ̎�ڂRK~f���;��s�a-d�y|3ל1�S���{�^�z0WΔm|\h�г��p���!��Wpat�P�ӭ�����~�][$������Hf�]�θ�M�-�}�Cw�J��e�;Uk��j�e(�
#�����Fm̧@c����=|�5ՙ�X��n�^���Zs:�W������jk3��ݷNp���~�f�<��5%X����a3�6�-�O������_��������I�f'-�a�r�j��a�B�x(Ե�5�~�'�Na��aG�6L<�M�N�O�{b�`VY���@�郟�V|���/�pѥ(�P6ђ����9������`R	T��/��स#��q�Z�B���9����ONp�^�O؈f����@�j�3{��HE-iL"!S�̫l�bס}�V6��3�ڮ��Sm:�VK�0�a.������<nI���M�Ӓ�f����sz.�����'U�y=�$-�� T:�.|0:qwbMN���Î�4��������y�g/X��������)����S> �@�.*p1�Z��C�%}�\I���Ѽ���;u{|e�U�ǶyÞ&u���)����F�m�IQ`�J1G� ����-�=?pK1���❮
K,)Ӂ�Vף	���������VR>�Z��n���mK�C:�g���}*ըz��9�@��̏Ef0��1_��1�j�.V���{�U�Ǫ{'�~V�nt��]���-� 5��ݒcm:s������~V�}3���f�؍�<y����Dy4�B9T|��Ҽ����69qOu:}�c*������G#P�9dRv�z�W�
jLY�$�6�RRR�?-_<�8���<��Ԍ��M)��o�K��l�N0�GtW��[`ќ�7�<*�"Bt�}�_��=��I;h�����Zlnd�@��	��r+*�د5���V_V7,a�>�^u0 ~Ճ�;^���e�]�q���������gϦW`��^�'�J!�Q��Q��UBV���&еD�r�P�����<'=~����cS�n�E�]h����C����B̊I^�P��[n��x�p\�b_�
��kcz|q���`O���X��e��E���E�iRw�U�}
7�5��Eu�é�n���0d�^�g�{G���-4�;!%̈́؞,2V�J���N&iPv�'�扥 �HD'��J�������){��W<��^��f�L����@�m?�1^�9:�~�����I6�;�\ai3o;//�k�,4�	���_֮��q�5���!66H�)�e��}۹�&N�^ڐ��_�u-���"�� #k����tß����,��醡�l�{O��}-�W�\��%�H���qk��À��Ο:���fB�ą����� �v�=3M軎/]/j�G��95r���t?%��{`�/c��&i����Ssc[,�(�k�%��؄�����MD 	���LL�9����q��]���������m3t�_.�[�j.�,B�X�Ł�����N�s��׼�y�)ׂ���E��Q�V�Թ_�=���&�r�fZb��Q:Z�� s��e;� �Ju���RPz�<��=r�ֆ���s�w?����-8�����Z�M�?e�����RdU��-�~ߣ�gs	(��t!��=g!�V��%SY�G3,=|�6X�>{��dSn�D��WNO��8�|g���qO�j��
UK
K\���V��G�q#�F_ �ߞЫ�4�
���{�*]�(�'�Rz�gqW���w��o��-�̉
�$�op��jp�%l�E*ްx�Er�\�=�J��"�����3��=B�F:�ʠ��粺��b��B'Zo��6�Q��{��.��%�	<mLZ��)w�@�_j~�P��W�l�Ѓ:Zq�+���.X�=�)��\�4O�ŋ�C�w/�4��,�y��j�7�M��.��>�x(y�e���o�	y�֛	GL:bt�s-����eM�Ġ�.�*p
�&g�	�h󳙶�{�ܠU�N�����7o��݇�����jOW�1��J�Kx/�����o�Ÿ"T$���Q`�C�`�̘���-j�%�`z��P�y�$�� t3��]ʜa����}�RT�E��2#C�Z���Z���˪s�ථN�:�(�~�,.s^or��o���_A$�z���+�S�N�����|�6Ƹ�� �]�zx/`�
�~����1iU5=�+����\��vbzS�_��a��f��ʠu%�8��ӏ~L��y[����9��z����I����)_��v�:������}�a��!�b��P�Gk�ބ$��ţ����%����
��f����b��w=NVa�2��Ȼ�9��v�ѵ ��ng%�r*��ղf��2k��/Dܷ̬���F��|&�ِa�B�n�}���\��8ƪ}����m3J�K�,�
T�<���Rv�K�e]&hS�_&Y��ś^r4+�{�B���?zХ���7ƅ�Z�B�P�n�f3/�1��b?>���P;h�2QY^�]�4rϱh��7�)�S3�v��<Bew���sm���S4�|�f�Vv	�^Z�ؽ�}�����5�~�_yݺ��la��)�D?�WD���9��l:��Mp����B�%���yA0ى��~�`��дV��A��a?9�C����8�I��҇섩��O�'ߺ\�|A�h	�g�ig�O'n��\��k��U�-�{O����Ll._ֈ$� �����n`�\c��^�`�_	��;K�Z�%�*4�B��+�FH��'�z9Ga7�T�e�J` �:9[��*�^��%<5�S��(���3k>$1{Rl$<˻�[�m���<�{�E��sdU쎱:�T�&5ڭ��c�s���9��;�p'��	�~O����#V�+���h��@qm��K�����8�̻�3�`B�{��%UG!�F�Ėee����^�~ס����N,�H����͒���/�,eLx�%�[蓼謚f��D�^�ƿ)�G��i�dϙ����E�y@��ʅ;XI�V�wj)�jc��ⷊ�����d����s�tuuݡ.my3�b�D��Nm�Z8�Y����}5+��x�;6q��q�|L���(�+Wg����+�/q��p��d�}�鐥�a��p��Q���WT�����*}~�i$f����)�J�8X�DҦ��mu�[�{1x5�$�y'6���{y��V������&�H��I��u[�=r+_����wfn�4��4�&��v��S��H|"��bf�l�b��9c���-��0�����÷T#�>�[�ʯv�6��亁�Hω�S1߽w���]}b����B��8�X&M�JG;2��5���c��������q��h�g�I����>6�j�fէ&\ �A>g%�O�R��>p�ǸV�HY�`����̶'̣��;��0p�#;׊�B���{;�X��f�E:�ٽ_v��ǩ�̃�M��_�yR̀1v��x>ܶ%�J�I �G��I��ۙR���N��.�"؏��h��ef��>Q���$�l.o�\`�3ٟE�|+K�nY@~ǚ��}��=;�����>�$�8H��.����~	'��ej���Xj>��~����x��{�\��;@�^�k���=�7��T����.�p��3M���N|�AR��LT\�54�
s�]�C��e���(+��%4�F���m��:|�(���Ѻ��;����n�����ϒ��4��|%�)������ϼ>�:.�h�㺲�ZͰs��3�j��������{��b��P�Зb�u�Ibo\F��(Ip���󺺄jv,*z"H᯽:�x�&��W���mB�EU�;����ݛ�"�SǦ�7K^��Cm��zw���Nx��Q��03lp��$��G[�1zn^VH�=���[F)�n�`q����qG�9������w_������c�n�v%��N4��Þ���w�3*9[�Gj�G�_���i����ι=�Q��5#��`ăe�}_q���� 7f�/�w<������k�r���>cC3�t�9���9�o��u���bϢ�1V]ahl�3�i3s9��N~�����){=�(⡮���#�~��*�a��F����M�G���Xt�Ø3�|�ǌzG�r�9X�͑��CN�܌�~�R	#�	R�xT�'@j�	������V��Չ���%�H���{ͥDB��8ߔ�1O���_~UZa�&��z���x�x
N��H��%���ܑ'���D(u{�b5�LV�a�����s��B٘E_�*]p.c�Ŗ�y��כr� %���]�<l�o]%�'��6`s����Z��#=��2A��>�e����L���B��@A5Ab?.Ϯ�2ĺ�b�P[�xs+'��R����MoIi�E�ͭ�C�/�'��@��		
��转��{z�P�o��,&l�;��W�s��0��-�3+II�A�L�H�����p+����"Y��]�����˙�q�T��h�.�>�{��F��������"�kk$�L[���$����>(�h4���gI�{ĝ�ȭrjh���ԡ�\
  �d%fbq�*���0VF}g�� q��J��n��I5X�o�&o�QC�A�0e����:����-pv�X4�uN�/l��� !�׃[�V��4G�R�g��r|��܅u���2�����Ȣc~�+`�牀P��_̉���WӞO��%���xe%ά{bV�X"F��&��%�wS�s��Ɔ����{�����pb��!��W�]'��}1�%Ѓ'�&aDBE�'��_�B�d�58�=��W|�M�G���0������x6���FHO����I�pUf�j�6�r��l,�Zq.���o	�X�y}��4��Xe5
i(A�A.f���$�Wbزm�[�J�ʤB��K��=��xȃ��w��;%!8]��qT������❯f��.�g}\��7�b��)w�4�^�}ї�>lh�
��R	V&�T �w�'gm&�4��Er�]�����ڻ��r�dh�f��D��a�y��uJ(<��z�Ո맶ȋM%#F�����xĨ܊��i����t��UB�� A����9�#���9���l	>��{h�����>��r�a���v���	g��� gg�{�/NS!oǇ�*��qY�$,݇,Hg!��U6)�kJD�na
%!W��C\wH>��ca�?��Nǂ���kz��� Ph9F��S^������c2�<y���(�-zm��q�6+O��Z�y{
]��G�j
�jD��'�ά�5~-�J'2�%2;�SQL��y*�.#��p��)qH��� ��bK�B޼g�\k�a@i .b�,�0�Nt�(�s��Dj� b(L��T�ʖ��y50����t��}#"��]�������1Vi?���4���D|rn�-��X�]FԊpE�x'ki3ڀ�fh�C�����(�W�埣��x۳�w�Ӄ:_��bC��sÁ����oRY��	)�4N�t��X-r�>ن���fP4[����E�Q����H}�7�&Xު�)��!�:k��,��KC�,�Hu	/����򀀌&� ��a�M��SY|m��y�ƮT����w�� �}J^�R�����Y����1�fΔI��K����M��œ}��d�.����ӫ��@,��Q֗�_C���b��w�a�o#siJ�i͂���S��'6h�ⱳ g7)���p�&/ ���`s
��<܎0w��c�p0h�h�5Qi_/̸�.N�v>��l��M�Y�1	�Q��u�/U�*���� �7ak�!x��E�wB\Ȅ���$TB�-?�8c�z=����ZD���B���A�+
~�Ϋ���`���
)�3'p�:�k����N��bݗ��u��}����KN:'Q� [��I��k۴�
�u������E|)Z��y+������"���W�q���6jl�7��=s�^H�ڠ#�r�T����B�{���:���H�z6tn���ED<dB�X����}ܹ���y���ku�bSP��.rE��_Z^5�G�x�̰��W	2����6i^!	�)[�(/�Ѹ���� t�t7�'�>��zIX��y5�[�uW��"��Wn��屁cw�C7�Q�7�%�~�������������� nA��g'�0�1�h�mS��3۷���.�A�N2l�՚�Fl��@f͎�W����8�u׺��q�f@��%�:���x\���d*}�o"�������SL���u��:9�­��:NL*C���ڮ;/������������[����B^����a�5�R	�.?���o|��^��b�$���h�m`a�*��H����PpX���ۦ�g���/�m���b<h(���B(�؆2x�輹^s<��u�'���ow)Tc2���;� ���I�y����K$��yEz��(�qY�5�11�oH�:�M��j�B��7�:�^��k+�g#ˇ)��,�b�Ȋ]��v�,~T�3��<��~��r�w���F\;��﫟�ܝ�1���!̫�S�J '���N��NO@��mZ�q��%r<�Oq(�&���fki<qdV�3�$C�V���5Ig���Y���Zu[�	ў���®rZ�wm���^�xe�����U�Ó�7��ԁn�)k�ѱ^؊y�vm�^1��)V\X��Es����)x�
RNcu7*��u����ő�'43I��b�ם2�}F��2W�y��@<�ic����>N��f�2Y]��Cz>B9��jP���bW�8��- H�D�
V��VS��G�[���~��s�/�����&�^��[�鈘���2��=�� Y_q��DY�Y���G6��Y���QM��9�(����'��9�xf/U� u�.�Rdk��m��k�R��,D&(���]�� H�[��s�
���O�__ �o����
�jxQ.��n�\��]z�s�@5�]t��ۉ����=�B�{���g5+:�<+�[�g�Z/���o�t�T��O�	S��Sǆ������j~K��G�W&[�.��q��#�^�ǩ|��OA�5�� �[G7�&�t�#�yW���Q"�/��{�0�龖���JS|d@F����4a%��|������zzA|q*D5wat{}~��?OωjA���-2h��6�� #�ɖ�׿��s�H��_�ϗ�g�B���/H�F�>'�I���$�i�@���7f�@��jED�~���"��1�qLX� ��R����~��<�7Wb�+� ٬u*��FLC)�?����r�� ���	E��x9��>�;f���a�\m?�$�a)����V�|�Ġ�C�/!��pC����X�B ��E�"��JQ>F��f3 ��cu�p%+~�2|p7`�J�ߜ��~a~�l��;�R�ul���6���	�{�D��[���|��-�Ue�rBAB�A����0خ�K1s��4$ ����@{�?= ��NŃ��~�'߃`���qa#X/tTJ��1aP*�JA�+b�m� B�	Tʪ��>O�[��_��S�<�b�Z������c�m��::���B�}`�ً�.1Pc�V��jd�b���$��|E� 1ټ]��J4ɺ�<4]�ܺ�	@
���@d�7�t�v�����^?O��tR�����ܔ��t����� 9Sxk*[h�����@6�ȣ%k�F���t���O����f�C#H��kSx6�����ܦ\�D�O�Ɲ�a��[�K^�D ��1$8��N��9�GZ�O��)��X�Y<b�V�ύz5�:�gb.j4�h�`�����`�d��"e�ɣX�7?�Y�D$A�CC�viN�2�n{B8�l����f��4���E*	h=���qQ�Z.�� �!'�w�/���F����~�Np���m�������"��w�_����╳*��*v�|=o_�=F#����0�a
8�4����i�K�é�1e^�4`�KxLj�so��K��J�ߖ��.���JǨ`�

��^fA�������7���-`�$� k�/�'�)�P� �bG��,��v-K��ϵ=ۄ(
o`�1q�GH�]����Gݔ�7�i˛\��
�
���GvE�s!jB����֤�v��ω�&�CL1�QH�F�_,d��e�΢�B���L�Kn�~ɐ��n�%��ZO	�9�)��]�S��r�J�n,E�J�@!�EI��	�h��K&�ԈY[^j7�ݛ��!��,s�4Qt3M�U*��:	�>dt��_��&����$-����셼2ߙK6i��6qk�h����\��_2n�Z3�<��+����'�Gh�����q���m�5)ȸv%y��$�Y�/-*�>��r;���N�K��zc�:�@Ǌg��&��ّ?ު�����7�f�*�fjܳ����y�璡�􏑙)!��h��l�AD2���k�w�&����1�/�P��aCd�� �@���<aG��	��?�9��B��>�ܢ�Ã[��a�9(�,���:P��9@��	��p�|�z͊76�҈$PD��>�B\�2:�w�ȵ��K���G�۞�!���_i5wRYԣ�m ŭ����o�B_l�5]�Ԑ� �&��m��3=�!VZ�cE�����ѓ�b�B�Y���${]#�w���"�e����F
K���JVPƺݴ2�an�J���1|ac
��0Y�H�H�����d�qx[%T5G�� sX[��[�*�(�hi��k[�;D�as��m�
M�j����?'��a"(�@�mTҘQ<�.��<;f4�g'?B������	'X	��!��Q� �4&�)(�O����٘c���!��*eJ�%��dkt#Y4}6�H+-qҺ��f��Ǟ~K4Uq0:���=�GrZ&C\Ȯ���K����u8	Zˮ���m�I�IU0$�N�^>\��aYrd��"6F���[�����9����ԛD{˟н�KcX���~�D��78{;�3�Q�&3_��0�w��cS�Q�Ĩ$^H�!�s0��%<�K����
�j.5���c�'����+��~����g�W*��o��,Eyq�@B����/�_I�Ӫ�i�g��c�����?l#ϐ&͈��뜕5fN���M�\�t;��z�E�ZrQ$�� *�؁�e��(�#�l�,Y��z��=^��4y�����3д�%�ޏE���8�"�I%6��}VQ�9�'_xh�� yD�Լ��O������d%<�:��Ơ�~��ď""u��X���*������>�DYW�GN�$
f����	�ec���;.v'��㺽����D��Р�A/t�W��&�M�#@�"R4FN����2�0�ra�p�j���Ѳ�I��0ʺ> k�;[ք��+0r�FT%(�v�-���;�q�AQ�� �!+�8*�"�6yj��:1&�K�,Bpq���J�FBM�o���δo���@p�1��i���<���DSB|L��8LR"�ABw��~]�J�vh��r�,�խ'���G�QQ��Y�%P�
����k��1��Z��"Q	�Nz>�.q���3FJ
ja2���B�(ѣ�=�$��s�0`di��pm���2��+����Y����2s�J˓vmH����U�aRR0L�Ӑ�Z;<}*�����^�ƍ�1�Uо��J�c�2H����F�Qc�|��} *~�P	%��Kt"5�+��I?�(�SP�0|�]q�>2j���&�|�!.w�� T
��B׷ �Ȅ	�S����"1�9����,3��{��>��	� �S��Mi�1�� L���7��5)P[M���9Gy�a{�B��¬Jh��Sy~�8+�͉-����>�@�!a�7#��[�0w�(��O%+�h<�)ƹ��ɠ2�mO�����v�(#��ݘ�?0m�+��|2c�dpt�y)�&�!H,�s �7@�hbz�¤��t�BF/Ch��F��po�����K�.o͎��I�_��p�BE4Nq���q������A9m?���H3����l��?%r��o�*J+N�*J�{�O�8��R�Z6�"	��͢�$G����d���+�kg�
\�
L�n���Fx`xt��+��ݯ�~��u�N>�.3hm�)�CY�M>O�]^�> ��r�)@�;,͗X�2ǡ*�Ƴ˸����rf
�&襳ן�����%+�˞�:k� �4�y����Z;�b�Ve�����sT���Ul��D�<E֑��M��1�_[[{\.��Y�'v�$
a,h�5#��5!�{q�dn�{c:�]V���i�|3�(AE�R9X6��ƀ��"Θ��6 -W�D�����%Խ�ݭ
�W��ȡD�"���KA����[�K����U#�/Ն��+��^��re���#d���ö�m��2����4�_6��_���
��Yp�{���	<��������Q�p3��������qF���9� ��k�:���y%�J��#`�:( l�'p��R��P���<��^�M��UK-t8d��C�����_DO�6�5-2!k�����p��0)5R�y�M|�hCu/Z��R��0*Gv���H�ly	C�3z�b��A	o�<�a� G�:�u�b��]��P`^��񋅚��%5G�9��?,� ��tD���mb|QvN�&J�p���:�5��I]Y:`�8�;�O��w_.�p/o�h;�:x�*s�U�^G�l�p���I<dd�?+���Z�x�mG}���;\۹����v�X>�׾/�k����@0��6F�m��g�/��u�mϼ����Ȳٲd�{�R��;�Y�@�M�$[�~� )
�<:,�d�d�<����^̀T�$�"��{�,D�,<�ijv���(cRm��3Ε5�H�fƔ�L��O8'����Z���S��rc�E�ͷ]��H5ܴj����F�mMހ+�Q���23�5�������'ohʆ�RP�6(�E	gB��B���M�s 4qH�T�`�D0`L�>	�
��IG B~���Qc�!@�v7 �
����!vb���_X��:M��w�����Z�4c��/QM�Wj =��ư�jA9U_f�@9Cy���I+���P`����|hc>(I$��Yoo�΀�l�x���I4� �싸a'~ȝ��'C$)<�Vѓ��%3W)^�i��b:�O��_i6���)���}p�Ņ|R���
oX��-���ޚgH��� ��pE�J��D�Y�@p�ƕ)�Q�XENl�h����rH�`k�5bR��9-E� Ր C2�8������/X�C��]L�
�PqF餝���k9ׁ{{��>Xα?{�׼��N��$>��� �Uz�+㯞b��Z���#+��]c�ˆ[�2��y��?;]����=4��ǯ���lIcS���?u�y���{��)x��S9F��ո�	���,9�^���`M�
 4_G�DLݴb�Ǌ�>�B�ۄ-GfyۇZQX�!J�B�Br��~�$�TF'�e��<\�p�T�7�<��%�y����0��J�tz�$��
�+?S/*x�f��ş�%�b�8CZz��;\:/7�Ql���]�X��l<��0��;q1��@X���f��Ƅy���X�f��1�'k���yXBm�6Qi+����#�Z�
���T������\Ï�~�8�*Ĉ�<���K�s���.̟vI��l���2=D���
Ka���V/�4�*/C�SgoT����7Q�C�]�;�ø��l�o�~*Xf�	�G�/���=�:��7��R�o��a�Q:��mc�x��f�'֪ż�����3H��Cu0��l�J��~9��A0�M���t�$z3�gG�P�(�� �ܻ�^��`:G���nژ7+k4���L��	�b{KT�j�F�� ,������ߥ	˫u%��Cy����:��Ǎ��'�c���c9eS.���	�?D����@�8X)(��R�,Ov��N���f�<0��
e�������F"�z{��Yp�>�F�H�������:b��5^�u�S����1.��!ڢ��G!a�9�B���N��A���j��&s��p�kM��X%x2K�ӯb*��W]P�c���d�� 3+��ε���u��8`��ວx[����b`�!DHQ�,=(����j+�6��������/o4���btF[�6�dm��
?9B >i#��;����|�psם�<~��Y�t��C�A�=B�o��/	j^�I��j�yN@�
zr�$U]���{�a���Rm���h�6���^�wϥ#�]�ؾ���@{=�=:$AA�q�'���(s��W�u�%8ǽD�1{��_�fl��9I��҈"�M�����jъ��6�p���{ n�[��h1"�z��$���67q�AU2\=m��(��,\q�����r�e���ܸ`]�-i+	�9u5$p�^'��9Ӣ�������ӡm��F�6t����v-���o�_�惇�����\�u@������m�D����W[�"�yد���{B��$�������mO%��l7�VW����BG"E�ΨCv{�h`Q���4_��wx����w����]�0�Ed�����M�oS[�%.j,�\.V=�8tz޷��k���*/����m3 8!��a` �xrN%n>�������R2�d"=�L}:ZGV� ��I�+����|�1S���O� �O��5N�|���r+tnFM�U}�:oPR�3Ћi���R���z!^������NWomh�����"D��(ԌKx����Gg�'đ����t�dH�F ��=�������״uk���J}��u6��Gb	ĕ�5���!�j�c���}��䶽[���fΞܭ��S���wG7O�(Θ�^4��m���	W	�ɭB��Cf�	�F���*j��";��ѻ
�������+y���sHF�kśH��xF(�Xh7b�^V?���-c��<Ʋ�9n�9��I��@���YO�1v/<��hQw����)��А�}���;|4>ɜA�������!'C-�9ݺh�7�O��j[�R�Mer�r{T���Φ@�M��Pi� A"'j��֝�f��F��k��I�;0HH-���%���O��*�04G����Ī:C���,E�34����y�.�0���ݦj�N����e8�3ނ��_i�UZ��V����7����A����2+p$)�H��v�S�����{�̸�[�U^w���^��yN�"e�m�áM�밦T�	� ������J��������pf�p|:�W9>�-�6��4n`�L �ޭ�$����'�1�L�)�8�un0Xނ�2Icⅱ���xLA���YA�zش���`�Ҹ-���߲���u�CV��SYcJ�����/h[�v|�n�4�1i2J��*��"/]�y�'<�qQb���ٵ�ZT�@M��G���&�}΍<7�sW���5M����']��{�>�U�E����n[�^j-��t��o�v�ww蔕X�\��_h�]�L�vⲾ�t�;�~,C|��b��=�qb��h̾�2&%�HD��9Lgc7A��Ch2�f�c?ݪ����dԸ�}�Fʄ��*A}��wIO�c��-Ěf�8�o�3I)��ʎ�(]��?o�5��+�~K[�Cx ���!n�h#^=Gu�����>s�n��I晃7`�!�]�$�{� Q��{���s�����t]=��A�P��?wZ�v:p��^نn,�����'���=����f��e��_/���#�F����^�C{!��6�6�۸%�^<n�l��aTv8��F!����}x�hva,��ЦZv�0�����ZK�*V���{&q��=k�b�?z<�����Yo��E�.��n�5��C �wwwwwwww��	�Npw�[~���{U�j�jwg����{�=�g��?�M��(0yK�1�Lv��*u��E6h��MuT�7�*Ȯ�|ȕ�Dl\�G���.w2���-S�q� ~Z����|Lgs��n�ŷ�:k/��G�{�6�	m݃�Kqs��K��I����$�O�l!�B#-��ă�j�y�bP_�a��.��K,��d/l�2��6�9�Qa�㉜��U���/h����l@�%�=*ZK��1W��V�ċ��2�����xE|5��<���)�-�\���=1��}���M�9���k�c���E)�7�V�U����N�9��Ӻ�_�l}H14�5�7�MU�=�8m� -�T�\�J�R�-tA�^�\-��%��..�/i$k�7[-��<�Q�
=�2G�8�����+�>�?�{|��(_l��xU�辆LR���W�����T���@�׏�X��0^��lg.x�����o[jp%uH��!��x$�S��1z�p>��ce�ٌ�k�`�B[r�8��Ka�6kFuD�����.��
e�*E˟TK�#l�D�[����R��Ƒr.� ��Qbv��*Q��P~@��>�d#��yj�~a!7���&�wܵ"�q�m�ڮ:Hg������N���m��'l��V���G#��%dR�呈�㠟�b8��`�̠�Z������Έ�9q�ݎeJX�Q�&�u����au�#t �>�P�ݫ�G�����ި�Hu�N��܄�]<�X�ӄ#�d�ڋ�����o�yL1�S�@Q`r=�3;,rH8!�� 8�,�ُ5�٬��}S���4�,u��^�]A%��<�x�캺N��x_���V����~S3�=X4�`�j{����'sm����m_1��H�UB��Բ]v)Q"��6���3rLr_��p[��p��������BK!�&�K�����wخ�Ko�ٜ���FW��(���"�b�s5�-֢�S��pc����r�r.���ɯzX�2���#��j��d���M#���"H�#��U�Fh�H�ZkJ�_��ߐ��c?�Q�;M��=�y����>"D>�y�� Q:J&�F�y`o uf�L������~>�~��Q 0����͎�_�+����bP�C6JI����T�q���n����u��q�m��j/�?��l5��	��H���a�z�)�q�Rf���iR/j1b�#��/�ׯ����C!��f}��4'��亵;���^d�/��%�X),8,����Z{f��IL���)�����Y���.r��[o�����>'1'&�0y�>���ꕍS<,���?�B�VyJXIe����U�`%69K���t���b�PluUsD�����	1!:���I��� ����_s�;m�3q���X��,"T_�.->`��^�v'���.��Vq������y@��y�0B�e%�A���X45&����iV~�g^R��WZ���t8),��$Ðӷ0ҽo~D�6"�����O�-q7LƓl�;��?f�c�ٝ�[]��[U%�W%y��U�� ��<{�V�ǣ�/J�!���.���|#����kp�rON�}��"3U�#�Ms���|�G�r%��\���	���Y����^P�G�%���y�|Ք/v_:��im���{�iV4].vZ˒_���yc�
�D�Zz3e�`�vY"�bʣ��9JB�E�<�H^�F��k����F��)�@E��]jf��(�+��58�'��'g�R��������Wヂ��?Fz.X-C���N�O�f�h�X��H��DS�y>��hbv?��8��2���g�i�o���)ے{�B5���ds�8 ���)�8b�\�U��|��a�J��7#\�I���C�1.@ߗi�M�뾬A�Y�׉�$�d˟�zܪ�Hߦ
EJ�rIa��J���b䎦�J��a �F��Z�ʪ�-�)d��5�(�W��JQ�P�͆���uC"���G!���{��E�f ��� v���X����і��8vU�m�u�Ʉ�󴡜�)���ΰ�Fm{BC��ܿ�e�?��%bSa���;��;r�ГqU8�� �2Վq$i%��qj0�<�@-5!��}��!�H��U,ۛ#�A�/ʛ�n1=.*����]��.�R�ٕ��H�v�@��b���#��� �����'v �%PCLk":O.�_�7!M�p
�(�h�s*��eH����p��Xi���D� �(�h��E������[R��=c���%�oPzb���b�9�K��L�d�-=�^����b��@E���T�ͨ������K������24�M��
-ǝ�,����o�B�.y�Kvv��8F!I���;�1���{��q�.�+��z��oBZg~���*\�ď��V�76�X3���#�צ�[���Y)+��"�Y�(̎����_�Q�u.��Q�b�:59�jM:f���#����0�����J_*
�xK� �$�`Ie�Qq����yV���f�"�#�0�b�#X���_���n���y�k�O��	�v]�V-��j�S�rf3`��R�ԚY �耱��BN\FR�D@ӎV��]V������ËVR�+�Wa#�Z�W�����v�
�g�3�Mi��%e�'� ��Pm��M���ۥ��������F�I_pI��~�evX�4x���I�ƾ��oK<�F8��Ҵ���������~�feb�
�0�s�I�Q"�}�x����e��T�'�wZ���~,����u��l}oh�>v��������2�bñ�G��{�acMu����ULw*z%l��bsd��� s4��7���ƥ�q�ُ�&�[{���^%-����������^��s�n/���.�$��b��%lG�?)sOh�*4�M|�N��#�KXJ\�8X�0��5��Ѕ=�{�]���"��nfJ4��� ��L�(��#D��9Hug���@(���jׯ녔�#q��v��HhM9n`i�����n����Oi�n�w��'ʛa�}3n��N" M(��3��6�L� =�P��9���n��n{�?�7�Ȓ�e�C���c���i���E:b���)�[�m[qVE�����cjd7�G4��?g�v����u��g�E�ƔV�A���>0���oT�=�_��|bc��@���&�ѹÍ)"N������7S�n:�;��M�ͯ�mndpWt�h���]f]�����
2�?W�^g��øT1V��τj��;��Hn
��Z�P�&��ݦ3�p�8��t2�5��M�haޅu�Rj��5Hy���.��^������h/��Q<�<��\�ԓ�D~�La�N�F�� �������vmK%����-mȞ�ŷ����8��^��GN�2ρO�2wV�O�4�qFH!]^�
@�83�@)�G8��8�K�9�̦��s�ӓc,�_h
Y&���P�=L���um�ZQ�lo79��|I�||!�QZ�T�9�,4�5јVl|��T�y&I=��|1k�%�ل0S�"c��~�+Ľ����|]@��+�N�ã�~�ӄh'����	{/�.���|tĎ<zJ��J�m^�R=���e�Q���z�fg�Bգ�:l���X@-��JP�t.�*>�8�����}��K�D�0�,m_��"����l ���9?|�'�9)�%.R?���˙�W0�P2 cb�%�dm0b��9�l���O��@�,L��%4Ɏ���J����\7�E�=(`v���lP��Wu�2�S�Y�Ğ�lֵ�8���:x�z������*��S<� ڱ��agb���Jv8��s��4��Q���6?"d].���F�����С�|�[�)��H ����r�����2D�>�FѰ���KU^��I��h_QRE�9oO��8:o�*l��ͭ�-.�w���9c@����RL,��.d��$h��J�X�na8�1�Z�9v0�^ى�?�T�;F[jc�l�i0q	��(4�3����ߣӸ}�J�y1>���W��.�����	�#^�����똉J5����&�4`���~�e<@[5PE:�	�^ǫ�~ŕ�c�?E���p'T����_Z�t�@��5(e�٬��JW�1pg���%�G�}h�-U�X���af��q�b���<�-���[�=$�
�,�����+��+�a��q��ޏ�g�;	�;&��d�_p�4tx���F���2ܘ]ʫL����}�wN�<Ԋ�]t6[y��Ȑ��9R>`�����7��H�d-����T6TǀҾ`�&�����|UKsy�7}�I�7����Y|5�{��9a�x�p���*ineu���׶1������#jT�������*~7~j���t>I���� Q��j���7��ō9J�u>"D
͇����0��� W����[*��߈B�+ ΢�hDx|��h�b/ڑH:�� �nCC( ]���8_A:sGH���q���X���l�Xo�����n�&�m��iL��ٺ1��'-"`.,�c!���D�w�����J�����D��ZE���(��N�*��Ǡ�,)GE��}��{/@�/x�\u��,-b�0�G��_�+�%��]�\7��a,<��e\�-�n����խ���o@�����J�滋H�"�	JD�M2��s��Jx��t�а�]�����$a����-֚R2ʲ��Ώm��i���-p�Y����O��24k���T)�5�U��L�^��-����E[/�W�&��T~�xI]�p7)Y�GBѲ(�o��)�I���^;U�[<��7���P�V?�Ŋ��%�i&�թ���Q��L[��d'���؜|�3�&�=�*�XMp�?;J�Mz�x�m�2��(cuz�جG#�@��f�R�\�%�қ+���-!��[��0�֎�y=y�j�=����>�;y|�v+���-v��{i9���j(�v9Trs�->v���V��q$�\���l�s1����IǇv��0s+�ϮW��S��R^�(Ix��L��m~㟹�%Ć�q�GH'�|0�6O�.��>�e%w
f2�*��K�X*��̮D,Q}��~V�5�����'��2TR���v!J��w�������7:�'=!e^�>^!}|�{�9W����JMa?nJS���P���1�l�s����wKo��UZG�G�=����\[l.-�7��M�q�e�xjj�o� �CiV҄<7�����ќ�K�,Z4K��K�ݶ���ވ�:Z�oNbS�^��#��-[q"�N<i�!b�UQ$���\c�۟�Cs�W!x(��G��U�)a2v��5�cԊ�c�6�I� O9�\�]�QEk��2'.�|��u��wP6a$ƅ8�EH�|^�f���_�g'���ie-��FTWĶ�_��Q��Ir;#�;1�~{A�6)H��%���/�bb9Iϙc�W��1_m*W0��a�&��t��S����Ҭ.C�6��)��oQ��+`�CDp�Np�c��̘�3�tI�gO\}�����q�{��l�]V����%sb��t04�X,
�&�,��ف�/&�i��e �f\�1"sЖ�Z��*l��-[��[�a���E���:�] gr'P��7":VD����?'��;c7<?�k��H�z����iP�J�(u+w.�5�w�6|���@��S_]���	�~�^�o���Ϛv#�kxk������%��A���ҳ�X�ɉ�kK�uGE0�U��~ǧIߚk�tU경����hh�l�a���B��sM�s�rp�e����� ����	D6�;|�yt�l�X��9�ǃ�dT��H1
Tk���F��m��	#{b�#�E9L�a���'����D�:��S,9קϱv�$K�|�V�q !�J�sN��S��%aD)!� B$-�|c�f�'��"x����d�y�\���#Y�����&{�*ӓi���wֆ��\��p	1,��Ѩ~��*n���ЛX�i��[��<ZD��g��iU�-��V�n�Z((Q�A�I�ۦ)i��Sk�N u�F�L�1���
��Tl��i{�|������Y!�;�7)��ӱҳ��4�S�(�+M�Nm-��*��_!�r�z�B�[y�C�2�\��{�#nM�qIv�1	��c����V��b�W�h�&�H-O⤯�3�N����d�PA����+��g���'</������B�P$-�̼�`�[B�0f~O�z�X��;=vKs���k��&�������A֕��*߻�;3�࿺?B�q:���i3��;)@�S�(��쀌�I%҉CE-W/U�����9L�=�'��pY-�����X�uQ$ѩU���E/�DQq�fW�M�m>b���)Jmgs?@��A-�o��
���l�j*�*]>�$eǂlu�ٵ��5�Z�e�n� �"����+{9F!��1g�{�F��
U��`��)�'��%M��#\�sk`�SĮ��}3���1{��&�^�`'y�J^MY��?
$G
�$�'�"b���ha��o�}=W���`�/޸�ӟ<Ae���me�����x$��h	h}m�\�z�;���u�nBCs��9�ޜ�6nU��)8U?�,f݋%���I����Q�8�y$�"i`�^ұ0��뚧^������Wpc�l��5#�&�6B���fղps���qpi�Y��pv���um	�MRF�*P��#�,!��L��GD �	�2�X��e��������o��"�_��J.��Ԓ�d9�I����B!4��qw;����o��ar��($�ĥ���LG��f��UJ�L��E���f�c��,���YrtZڮ_����F��^���B�)pw^�w��}G,:��PC�����m�P�rY�_:�%��*�Tz��e���R1
�R&�c&#�&
Pj7J|�=�,�ӛ����Xy��)3Hb�7d-߽JĹ:�ut��D���4��~��w3��[浻���3�$��bY�ܟ���H*�y���cdKS0~c��@v3��Z��d0p@`g�p�c�#qDSB;����Jk���K������ލĪIO��+�[��M�����E�=5]L�qO�f����v&���,��\&�����&^��"wk_�6/�����'��ݕWh����F�9ոq��qL�+���ܨy�ti���]�ᢐ�ow�2Q�}���t�襏�T�,��ދ"rz���g��{���B�΃�+C�5�,y���k0@0$.
��b�;�laS�M��//�|S]��&V���-�\	�
Ib��Q���"�wg|��x�z���H�w�Υ��;��KiN����������	��-���?���\,�č"j{sS-͝{���һc��q�� �)f��']��-g����(�O ��S/�f$»S,g	������FN���j���u���9W�7� �=hHͤǯ���m�� p�}���`B��W�'����b�t�_>�_�D!�Q����4��νkzI-�L��#�Z~�;)���q�
=��P���%N~R�3J�MU��٦��`q����j�<`
�M&�ȃD���Sk����"q���f���i��tv���s�(0ahG�,����1/�[�����:R�"�-�ʢזk/M�k�߸�ܭ�G�M���+O�3���$�zЕ�{a0�+9E�ύ%B>�~���..�B�%`/:A���M��+O��[5~�[�3��_�����BvOe��e��K"�"m��D⿳甏����5j��g�yƆbu{�����Z�X�=�X$}\�.�SQ-�����/7E���豨5�Y�%g`<�~�y��y��_"�k�P�<�@�p{<�'�m��(�����T��m؈!*6��1�s��U�Gߑ�{�������W�	�qDTf�,�eu�@�f�������R\�{<l�1�<�W}FN@N���D;x��b
���vޘ@#�֞G�s��p%��B�׏�uW7��B�����*�ƭ��KC�zeGТ�Ұ���۩�\�A�E&�)_2C0dKj�3��<��*Mʛ�2ul����gJ&��b���o��֩��:�.x��!rq��:?�+��ä��\̔��ܯvɒN]��Lǝ����9Y  Z1Ls*2�m�)�J�{7�|����~����f#��A}�������nh葅*:<�Q<�g����3��j�v�0�ߞ���_-o������t1��P5fW�Q#08�y�ں�����'�����b%|�dz���-]���A��ҳSgɪ���x��G����]�=��>#�n������z�Y�$�$f2jYؼdTk�j�Ȩۺ�>��H��Y�z}�'cv��S���Cbr�0c]��zb�c�S{}�Jq��R���8s~'�rg���z�_B�_&eϚ(�&����k�Z(�'�L���e�yND��r#sf"!���.9´�#������N�l�W��0�>j*Z̙��l���|$c��.��<	#�K�t�%�]�w�W��d6\���E�!h��cQ���+TǱ��J��)g*�AO#߫)@�F����#j��Dv��8�1�#�������
���������q ���C���{� �Ĝ���mT��N)�bN� � u��T$h�TA��!�O0�>;
m�l=�+9o��i	$ĺ���L�9X��]C���!#��U�Ow`���_��u�1I<B�G'h����j��ȇ����������;�y�/�c��M4����D���Wr-g���TOT��x�Wqɑ��	{O(A��a3�\�to���F�l�d�)`�/���9$�1Sy � mؾ4iYzѼ� 2�N-U ��v
�� ���O���w�G��O:,\��z�|���������=�U��W�K�?^�N�9��&���
̹��D%�.ѐ����-���r/��8��0R�e�����3�t=}98)�PY]tb�1��K�U���&�-F��:YAyg&���'�?_Y�[�C2-;:$K�J)~`�SN��8n���Mi	���%	cA�����
�y���?W�B�e>Uf�t�({�����d_�\ŬI+#+1;��fD6��Y�Vj#��Y�L,Cf��/YCoȃ��P�5�AJď���<a�X�����Ȭ���SN�L��z�1r��&�p�3d.dm�;�e�_z)���?���<�S�嗕�b�/^��A�geM�R$D����1�Ox�!��3�#pKv����aT&;��U�c)޿��8/�����%%�h��|�j�i"��@#����槟�ŭ�
	ꏜ�^{BHaRԸ��r�ɼ�{qq��hF��/r>��~���.��G��f�G���L�LYk1�qY��g�J�LS��u��P�!pL��_{�Ĺ�P�ٵx����nL�n#�z?��q�[/�Z���*�����"�c�����e�]�{�2�ȂPəE0����,5/ϲa��җڌ8U�L��6��W�2eM����pG�3#�5�|X��+���"O#DôZ��5��pk�(�0�e�����0��M&(j�J��䪟�k?�����dْ�ēz����~QT�͇�������P�]R)�;�P.�nν�ϻ.��Τ�{���0v���B����¦�m�a;#��T��=���͗�&+���ݷ���w�8Ʋ�<<מ��41+��+{)��z*~��ASJ2䍄KV���JJ��&m*�9�ЂT
8  U��ͩAEh|�e�Pj>����OW��9�T�}@�\��9,�t40ș�}g~�p�K��*hV�)�$)���>>��DC���E�@�x�gE��1�X��s���i�E��ؔ�6˻�Iv�l&��r�����& ���筇j�k5�Ъ':����-��o�P�g�����c���e:/;Cr<�#'����w�=��H��0�L�hJ�~ ~���Qo�)�Ջ؁����?oMtDx�1���g..�;G�z1�R*>x;�u}�>����歐"ah��[��x%@a����|�������(Ll ���/���1izI�!�4�:(���v0�h�����ï;wU��{�6|���{�Qq׫X�q��Z�m3M��1k������P[p>�����V'hP��(p5��Q���,�� %��+����&eg^��������L�Gw���X\
��)�q��r�O�$Vo�������'�4�7˂e_�ּ�_��2k��-�1"D\�)���
��X���aq+m�(��u+]���G1�*g[�k5W��^�������;X�ͭ\	I�@"d#Z��4��K3��
��Q���U./��Iw�e|z�eSl;\������x�:K���J~Td��>���r�uPuh��ד�_1�#�ƨ����kbJ���p���" ��t�PW���u*�&�I��4���E~z?'Kǉ+_>�߭x�P)R$b<� I�
Il�´]�������p�:�[���������PM9*a;����z�PRD��>�਀����=���p\��v���N^
LxLx,5�����G ?=?1��$SK� �ګ]��*F�l����ϊ����ˡ���]���������~9o!X���Je���-��M40ޑ��D~  �VLPL؊���WH��i�F��hX�O�=�K/ �A�%��Ȫz6^�R��q`0�bd��ۥ��x��b� ��Q���<�ta�N�qX���H<�E�-�t��L������F�J�}�<�0���%�v�8��v<ѩ�"��eZ���@C.O�������`6d�[�� ( .�����F��%��'ؒ����Y��cs�m#EH�/�^G��kik���ʡV�1HmZ2����k�����^9��x1�"�˺�~���V�Um��ڢfG�
�A��(�D�__B]�U��u� X/��������nb̌��H�T�P4�+Ѽɔ
�e����fz�-C�K��WSx�qh�儚��m��0�\#c�&:cZav���ƑL�eX��R�_8�Zk(�(�MŪ��6�#�q-��~�����	��Z���c�MA�y�E3����E�V,[��(s_Sf�ik�2�>��SA����cg���E���ݍIU4������e���\� ��_�Ѡ3��������%S��T<�(A��e�����rG����J����i��[f�v�0:�D�kE2���m�F�B�m�K� K����B�x��x��@�7�g���ŀh �2��πx�`9b�	3$3#!A�xi���Q�f�'�@r%����u�#Z�cƔSH�n�"����#{��O��CVB)=`d��H�U
���d�����&i�����W��F�Hhp���)}�+���B����9J�������Y�>z$�;���IH�(��tc���^ϊ(��k�A�[5��:�b��)������ ��mPI�g!����i�	� Ɓﭡuud7X����Q�Q6l���� &P0D��k�1Q�1�ݠ��#U���/��	W�4�~���|����������#0��]I}���~22�8ZN2��2#q��|�P9	��=
�H/����C]s���O��WD�;��B��f#�ϻy�ʳ�r?\�ӻx�y���&���pX�#���ٮl/�cW�O�?xF�֎�֮l�+I�+ǁ5l�~C��|׆�zX�jF�CՅ���?r�?��$�%��[%�ȋ@�zbB^�L�����(�$��͛ޢݪw�@�:߅��Txa�p�����p�a�XwJ�R�':��!����Sb����P�|h/n�?)�5Cd�,��Mb�ߠ}fŊ,�W���H�|+�0�^�:�;G������Waq�~�_��/4)��E���Ç�Aq��5+Uho33��$lt����S��|qFJ������9����[O�g
T}��8h��Q9�P�/Q!�Z�י,ĥ�߆��A���q��9��cbs��#U�h"���D�5�����季47i�Pf��ry�L��-���y��u�gcN ��R-��<2�����-+�K.
�������m�p48(��bwkw��/E
�b�+�p�tL����,uP�@�G}�LfE�"(ѽ��9dm�7;�s=�bD?�nD��f���6�L~j��n���{�׫᧸�.�uю�`�xΨ���`oE[$�����v�ؓ���r��^�ʙ����<ݩ�1X�ʐۇ�ё1��a��M�r�)��=�7���eOj�_�n�[qVcR���k�"�'RS͆^t�q���6������F5��Ϯ���z�X���f��l���e�f�:�>|<�?��{�|��k
 ]#�a9��F����GBKb+��h��L9��x��K�Cػ�������2�<8Ć��y��u�^�~�7���5q�@w�G�d����;o���oy�K.��1�}X��QTh��Jܲ���j�H�M���7���-$|��\>O]��(���ܽ�7�2;����y�<>(m�w��l�� &��X��V�$�"i�c��	��K�Pt8��5��5���"!s���Aqpb`�}r��;@���Y@����T�P��ϡ�j`[C�_R~�4aG܃���n$�/��������/U����W�߆=%�-�B>O]�����<ޠ0�[�.X$z�`���>�XXx�Do���0����sx��T����zO��f!�/�VoC�QZ'>��5�;��p�����٠3*L���Y�Oɛ�/h=�(b�GHl"0�,x�,�	$o7�AHm��,kM9Tcc'6*�V��Q����LM��u�X���t�p1��x��s���"�Q�k#��� tRI��.5=��D���"*�G���n�ϣ�DC2���WR�k%R9A"��w��

&TM�0���kZ�g�#Cm0<ZJ9�䢳�j� �:1����;���n��GJ톌�hS�	A��/�(i!Ԭj
Ʒ�XQ�n��y������\	�"rҐ�����U�l�@@�耔?�U���$�����?뚌K��,��7��#�<Ba�M���c�������	v�j��Bl�����������v%5<b=r�j����ك��3�Ա@�b������inQ"a#נ�a�$��.\_8b�n0��ē��+� ����"�Y&�
V
�n�x�]`��?-�@-b০ޭ௠�h��s�&Ip�?MP�YU��_�U�>�D�W�'�^[͸��J�7�� �\B�!�����48�9��̥�F�:f	t��vZ�]�o��q�a
������՚ax2����԰n}X���Y��^�A���&5�M�
�X�O=^5��ضN���*W� e�����4u��Ll����F����n�i���h������0[H�]	?G����@.j�Ttàı�+d��rO��� �c�-��OF�+�T��ϣ�9X�
3��Թ6J�軱�i&C�G�Eώݘ��g��I��\J+(�z5l�s¹3q���2S�b����ҹ;\���F5�:oF���&��0��!rWf��5��Ħ+J3� "�{��P���r�|�Ⱥ��B���yz��%���LF���o�`��M�T͢DE�zp%�
x��[~����$��i\f��1�ǖ!B+!|��_�(-��.a�O�~҂I'��Q+gWF[�ȉ8h���~��{��;-���9=ul���W��N�v+�>�z���*�R9AZ�=��x�'����*{�[��k�䷴�� �bu!sZUC-�a��g:p�:�+T������=�Q�v�B��@�S�t��R�ڄF��^橜�e(��݂)��1�����t׮qiΟUmڷX���=�Nz�$H�9t���1X�B�X>�P}�?��d\��	ʎy��xZA���1M�%��U)�ک�[�U섎�@gB�Y(d�7}�����[Hn��lPQ��2vvĘx��&�i��{+�X�"�'�����=2
�i�`�U,b�gf����G�l��"�#����xI�;��鈸��A�,5;@F����*�P�m��&���������V�k~��K�- ��p���x�n:�>t)� x��M3�)�M�l8�-����KG����8�`UI?���`s�F�p�2�}Z�����O�Kc�f�
�!pӪD%���׷�H�
�8}�Q/�`��>z;C���49fjEPo���X�Dr��;�5���^�[� A67�>X�R�ny�7i<��PI˞S��xMx��n�X�_��O4�d׽�0[Pr�eT��⽬�k3<nvGV�P�^.�/{5^�r[f̉�6�y��y��E�YE�G���*���Ur��%���`��Y
�Ʃ�@�����F1n5�}�z]��<.�W��D,J�d銛a݇�Toud���:D��Y�$��6�+i*$�C��`�S�ws�c'�]!L����qZ0<��Ȃ�u�Nw<�����D��Uo9�i��ş"R�!��,;�6�\(Ճ>�X�>�"\祫=�Ǿ2���`����_i��S̹�1� :#��j\�����[�'��f���ن�V㴴"veў135=���	����ɧ��� M��`���c�5|J��i���'E�)27�J�㯐$b�)��B&)U!���f��A�m�4�!b͆�qi��}�����J��9O���n�8��
�tF^PG���x�\�x�[c�v�RP"?SJы"��q�r����$��Y�l�(�-�P�J1��^	CM}h�T0��	�P�Cj]�P���C}a&��l���Rگh�����@H�.ޮ<ֹuSC�˻Y��h�Ш��R���.���=�C�X�;�J%V�ik�W���z�m�z1$ވФF^�7^�'ۂ�1����j�B�tJ`q~g!t )c!�B��|�-�k!�Q��O\�'��72L+�|��[9�VX�7ڤ]<e?K/��@/W�Z ���d_-Du?Z�s�S2�&:�#�$������tJCe��U��M��;��F��x�jdwv��ѐ�8��7�
�����1��9�-����"ɅR���48k�nն-��\d�p�=��zd)�hk����ۧ��+ �mT�v>�w�t��7=z�ʁ� H3���F�K�#L����@l�[Q�����6�2d<���'D�T�F���-mV+�#�&��0K�R���k	׬��P[f�_AnWL�ˑ�U*�u����$�zfz��F�Ah���B�Ǌ7x����ݰ"�ne��u5�B<7�++�����20ŎW�6�<����ܑuk�����\�@�B�)+���k���M���J�\KFg�"T�"�E� h%�#�T�  ����x�B�,\�b(g;���}]�@~ݍa��V���$��]�+9��FM.I���7��3Lp�e��sfn϶���bs�+������X�4�y��� ������8�����"�$�	f��ri�3������MǗ�W*����P��'R�t"V>�!H��.�҃e��8���ܳs1�� �뚋��k�6'}b̧���3�!.ko/DK�[Q#g7��e�
�E	�zzh~�p��7LP���-fv4��?�L������5��zw������Lӂv�~�F�:xe�~��;R�r��|<7Dת.c�~(r�h�r.� 1O�$� 3u�fj����(3m����N�>�l�|o�)]!�K�r��?�F�ڋM�~��u�������K�$��8A���F�ۂB����E����z���%:|���Tcnt�Ve��=�)[�p(���O>2�W���u�m��Nt�>>H����_C
�k�S������I�/��l�4B(������Q�lcNx���#S6A�s�d�m��6j�-�-,�C�7�Mr�x�61/x ��QPR�L�㱥��;�m��(=���
�#���ǥ%Q>���/|��O�,����F����\T��L���k~j���@�����u�.�"	������G���Qͭ��a��:��e���>�6���m�NU�1���a/�����d�-�p�ȟ�t$*x�hgl���{X��[7#�3K�*�~��Y��RN�7*+�	���J����L�������Ȏ�rO>x"�.[M_�	_���/��SD3���/�K�+Q)�РK]���ճʈ� S�K�gf�܀+�D�k�y8x���o@ݬ�	(����|�#� w�8
l>��������3
���f&����Z)�ϲ�"a��V�����' �=��e c�8����]������0�O�h��y�"�������W3M�A��\0)k�ET3�q�0���>ҳ�=FY~>�����:9�_t] �;�ne��O��/�X��R: ����uЛ�Б��ۨ
��na��y�&�{�RO�]��p�>��[
�R>�����I�d:�H�N�1�ż��՚ghM��h��_""���<��lHaoh�/RW�;%��Q���g�J�r�
�F6�1�9x�m�����+���0ww	��������5��;!�����n�/�n�{ﮮj�v�gG���z��y�?(訩P]�Se�[�P�x����8�>��R
e��c^MI��T���7�#�ʌt4���h�#U��NKv%�9L�U�.��9�U����6��V�B\�ِ��H��b��}����"y)��tϢ����m�[��^L~ng�p���;D��|�fYg�՚�Z; -<O2.���{�;�� >���Sr�$f�X�db�ߧ��sP4�AF(8EH�v�ӧ�%��&T*T�u㋐R�tI�=�����U�|L�f��]xL�.mL){Bh���$�-)�{���ǩ�M�++�M��d��G��ik����@%߬5B���Tk��#l��$
y��f� �����*~�~	�h�*=Y��fܢٴg���ǐy�Cذ�	gT�F������~*gC 54�C�/��$6���y3�^yG���>L��C_���W#2�#���8"�V����z��hm&7��sD����T� �e��Js�@��OC�ov�$t�)� ��*�@�Xտ�$�����%�Ù	`<g,Ql,�����S�2h�U�|���e��Z2]C;���s��N�7ҕc�~�Q:B�$C[���F�dn@L����X��/��;i����%��~l�*���L�G����k�
ޕ�F'�)�1cD�9'Ș���f$���F��ؤ�W�_�c�>oz�$񾅴�E��0�����*�7Su���G�]��3(�U
��'�@x�*-�^чY�ʎg�!�Rѹ|gCĞ8�̈ޣA�
����o�J�%�)~�R�x�%I/��̷�I1C<��20�kg��Ӵ�l��i�d��CM�3�_�D�<�|e��O�kII�_%�j�^7���L��ߐ7�T����B�є�D�C�|�`(����e�B��8�-���F�G>��2�E�	���K���C
�t���$C��;�5�uQ�!.rX�W}�҃�YU��8ԳZ�&�{��ږ��x�v�Nɬ�;S@�G�P���%���d���x�|g�}�t�a�OWC!�R���~V+�P����o�HkbX-\5��՘�H4�%e񵓥����~�����/nO�[f9�n���	�,	�x��r��Qgְ	�(�pH��$�5n�>(�}��'7Ϭ�{q~�솳Xı���!�\�����.$h>� X��S;ђ�o�~����a:��c��pzT��榳����\|U0L;���L�pK��%���s��.���v:k6�ٱ�R���T���3���Lsь���K�o�9�����s7�\~�C�f�*�h"m�QQFK1����V�u�0�,�#��Nvc}���xC�9P��C�_8����^�&<`L��E5�ٽ}�޾%�_zJ��dP�7��C�U{s�SP� -�e�l�hG��p�T-�Q��:��tw��d�f��j�\�"L�����'�е�d�з���J�P�B-�Y�Uh~-�� ?nrN\���8�u3�7�z�^jԷ?�_i�uJ�~ū�)�����nL�]����`�:`��|�թ��+�l����+��k��'�R�h.��;���**#�0��,�D���78�)��%F���EV�*����C5@����P]s���	I��Q���o�i!=�A3p�h��I���
e�߰R�y�oR���KF�^R���1�����y���� ۛ�I�(Π�W���8�#m)K����ۃ���x���=-������nS�8��ܟZ�&�D��4{d����;:?d�T��z�����k��I��Z�����an:��ԌP�����7�g�c�fE�5�[���M#G��D�<U�����S��0D��ԁw��+TDi���)6;CF��5y&Fzc	2�sr1R�p&�����鮆R60��T��s��\����|�~��������U��cs�ϝ�>]��ރ=.�i�g	���n�x_���BI�L���IoƔ�C�^������RVDY���ܞ�����5�^�
ˏT�|��5��T
�Ԃ���TTV��t�G�)���6>e�|g���	I8�Fm���S���^[�n2@��ݎ���R/O�+$��nn�-�@,	�����}���`n���4F߅Rw�� |�� ���X%�R~�T%nLO6	��4�df�w��[��,!�[Du��UŬn��!-�����u�N��ςz�m��\9����wh�`i���,�Ҁ[jz�3h�rLJ�0vۄ����[h�+��FE��}A{Rp;����~f<t��	��Qmk�Ty��	����ַ=��AcB�%�#�c�8
��?�m�v�	�N�VT�3��C��}��Yẜ} 
��(J 0�C$�V��+	\�w�%�'T����l<��m��G�#�Y�.#>a�X5��q$��E�����D���`�{+�#,��:yi�8�=)��嬿V޺~��m�������:b�E�$�*�Hۆw�Z)�n��t��� �p�!��q�B�"��椴�X�Bx/Sx#��4x���4������*�ɟ�`@;�$� �zU��M�(rtd
��u}��d��/�J�3Oy��T��s����l>|p*䣆j2E����"p�N$��H\h��F��?֯,ܘ��P���+R��*w�P%��o�I�i,׎��a�ƫ�������$	�����.�RǦ���>���,�D҄&���G��k���w #�
á|�6�µ� |R�._@ _�FV�>>W#/������_B>n�S���J*fk$p���|�K�j(��8�Xǖa�x��q��eG1}�3
�//I�:;��	\����8Zr�����rE/�t!@fu �^������?-�q�I�F��s
[~�����CS,&�����&�0fp���ٯz��H������=o�;��vgUř�WĂh�@�5q޻�0j�d`�O���ձu1����e�y��!��dZ��`~Ÿ����C'�MR�t`��#h�#.G����v����*?/�����^�
�N�^8��O�2������&��6d ��w�m�LK�c����pS��Z�ڨՌ+KP�`p���=�ТY ���1W��9V��?\�����\�R�\�V�s���-��av:}�*�����[�s9����EQ֏>�/�	?��f�̻[��	�!%MW��xm�d"�Q�SJ��� i(�A��~�Oo���#s�&A���|�ЁDϥs0>}��r!�*��D4˗5(W��|��W>�G�ợ4��f4/��e�s��l�I��H���]�t,ymo�~Տ�Nr��t�=�Z`n8�4���k�L��Y����������{vN8?�0�z"�G�W���`<����5���>�,.��(d[3B�:K �;E���`C��hO��,�$�J��"%���X��q��"�.v1���iP���Oc|�C���.�+�m�c��|ٰ`k��ƈ�k$�� tC�e6|nի��4L�'>�t�e�-�$z~���;���+�ֽ��Rm���ZZ�w ���JM`��&�Q��h@�U)%���yj��0�G��n��eo�~��m qE;C�;# ���/���B=�,"�
'@�%��G@{���:�J�:7��E��=���Ly��s�ߏ��\!�~sv����F@"թ���5���"�I�|����n)�&�ϡ���s��9Tb��OPվ�s��"s^�5�%�A����D��p�FY��O���Ѱ2�rI���h>������s���]o�TR�߽�u��z��������t���"��ڱ����?�p�a�fT���=�r�&Y�ݑ!����S�G���bw���k���(o��x
�d<�+&m�D�"�ȰPK�{��p��ѡ��M��S@�q}�=h�ׄ�y>L�����깴u����A*W����0K�M?�/ j��m��{T���>xVf}m���rh���\��\�U��pl�XE.�l�H6�Js_����>������8���iX6 -z�˴��n����MH7b�����7[8��M���K"�`����d is0I�hQ-����,؋�Z�:c�ݛbqk� ��{�|�����e�������M.s�����	��3�ϥ�� 	hW��9с ��k�=�|8����ȡ�X���Ĉ�s��wmQ�&R���[�^t��7��m�%�u>-iӌ��V?�`�����c���ܴ��x���OtZ�@n6ȁ��o���ra$����\|���)���s@����)����/�$�3�*	��f�9��uz��
����n(WG
0Fj}��[@<&���q��lq�L��[{I	�ޝ+���w<�����KK�Ʌʱ�ރ����E�7�ű�&	���%��-lHZ<����t������PX�mݤ�����d$D}K��5�%�+�L����Wk��mG� ���]�)��G������m��n6�L�f��[IX�}T	�]Hl��(S�����:=gư��I��۸�N�'��]�!e�pG=��Iq]����C��bܓ��U�����2����+m��{�`jq�h�FYv��Ajn.|��B�"0^�.�!;�<)��\3ˀ���.Kjr"�gCu�md;]i4m�?!/�ܾ�$��N7�X��1���CDOBM�8k�A�e2-6k��&�{˓��Om��My�ywvv�����H�|�)��TgF%�'��=k��=��ïA�`�KQ�ZT7q\2vk��U[�!��7O?��]"��a�n-��:�#R��������)�x0�3_f��
�D
��a��NoM����wx^���S1� �߲�.9��_��MK�v�aJ�x��d�
�,Y�X�ȫ��N�=�]�7E�3�E�l}J\MCV�#�b�>��=�CM7���c���t��A#/3W
����M0�[VP.�{����9�� ���Ck�O���h������OvEߘ�̷��&�I����E4WcY+���s��.7]>t<N@ J���g�z���Fce���)||�.��Q�5�,��*��$�C�v�Z 範g��d�ໂ�z�-Ԯ�#�a�T,�h�[�*K�P=��C<o����u��B,��	�N�����k��6�z8z�y�L�ʏ��ټ��S��('u������hؓJ�oع�ȅ!ӑ$�O��JM��P��!�Y3��Ƚ�3����ɟ{�,9�{��Z�����������d���:�Rˠ��%�e�bg��uD\𖾇��gf��8���
�[qI��d؜�P�.����4'H��P.�Q%|t?��"�w;��Ҽ5�D�l�&�Sh�J��Q��F��~L?�ȉm�s!�A��Z)�޹E��{ۇ�G���8������{���J�� ���E�#�������Rb+�4`L6�G�|��F�K?��r�g��IWйH^�q-Mn�s=u�۔�d���3�&P)�t����O������x����I�g%~6���Y=������5�9z1>b��O�G�w?Q�|�LP��l��U֢|��#Tc#N:#C�|�v�\>>�Dk�W_7�&P�+����^�>y�ݳ���W'�Dfh@5�³mнVe����[K��B�6���]���u�JJ�B�:9e�q7����/��3*�r���8��B�GjwP�G�U�)��ſ,��:W�;��qaݩ8`�������%WQp�])���Hʼ���G:� ���ViN��S�D+��b�6�?�a���3?]*�r>h��<��������݁nX��"r�*���Ɩ��˕|� Z�A o:�?�x����>2�~���l�#ξ3y(��3�V��� �Ԣ�
���7�Ᏹ̙8��L����徾��q�U�s>�p-�٥{,�˔x��g�Z���]բ���/���,���՝���qsu��`BHþ����5�[�ԅ�������|�A$�a6�$fB���Q���5�x;�F��G���c�B�
��6";ĺ���
��oW/h�3�x�K`����\c�Bם�ul�s�)﫠et���[�U䌄������&�܌n̯g���(`�E��rqqI%ѵ�n��G��$p������Ͷԩ�\ �e���R74990�؂;�+ֺ�����W�3h��էBO;/Jb��<��������[�j���刍3�cM���B���⺫�Z�|�s�7��}�[���Sjf!���sy��`\X�ɾ�~^�k�VeI;5�=R%���V �g�#Tk���C/��i��!KL6����ˤ�h-�)cv�5�g�QB9uz�>�0D4к������U����u�aA�ns�KE���Y-���:P�I];�����@���/t�=.�r�6�ʧlj/}�'_1�
���P��7� ���S�l�����r���$!d��tpXr"�Z]�]��^N�(@���9��t[�Qvz@��fD|���$����Q��{`Ne��k^l���`YJ�=s�%oqg����������៾��;��^s��ȥϴL;�e1L��(�1|��{���w9!n'h��'�]3h�]���
�
:NЋ������|�A��wd�(��T9�c�s��*�M�sd�����7�To�a�.Au���H�gZ <]��ĭqǍ���C+����廁ҷ?�ڪ���&�bp�)~��2�/ʸ��45�e�Ҩe�h����3߹�<O�`�F��ߑU��0Կ�z�q�I�ND��w�xq����PP4�d�n�]�<,���xI�:)I�ވt�|�o�7P��?H���cסMA�t%C*U&�m�����J�i�ONI���9�%�S�����y�H�֮v�IU����bEq'��<�"CKh�,��IM�<��NȆ�h1@p�8�D��t& tlg=<�X��ИKԡC��;���{p��!����Gڎ�������o������3��j+B�����۰�f3snbxU�|����3p���}�
ɓ%�I��n�N������M�&�8�ZP��eԸeذylKM��.B�"@���*'��M�
��=�CR��&�C��CY��5��M�n�
�.}� T�<!��s��(�G�f8�+���S�'e~���$�-j�yk4}s(�
��F�:���{�!ʫ+�D*6g����PTs1�5��l�uR�&O������d5�9�И�=rũɱg�)B���ir�{8#q�����3CX�{�f��M%�x`�'�BP� �K���lI�����9����_���9� SG�;���0O�<�z>�f� �]������D
�f+�����wEy�ǔ���-��'0��w���,�ʌ޿1�ډ�� ��d�	L��䧘],��|�'P����S)Q�;mTq�О�H��.�Y������Y�/�������� òu���j�b!P�4,�6c<ܩIs�6����x�ݹ1��ڎ��J�,� ��%���18t��E�&l�4<E����F�[�5^ٟmvf�2��˷p� � ���<��P靯���˸dG�>\w,�F������W�^E���Jx;��=���/&u�7u��r���A���|���ɼ�0��1���r4<�w����ƪ���YE����z��S}HYY �҈T��Z���/�:�E̰qI����:���h��;��OƗi��Y9t�w_ �|U����x�]�;�Q��<�?��<a�C�-����Ҟ���E�X�|Ę�{�rL����ƽ�����'��$v�I���l%!JU��G,F.�"�|P��i7<���G91�����-|Q��:�W����)`��2��ǔ������^�t�O+�X���xzY��1ҋ$�|ْ|�>3m��0����/��^��6	�(��V6A����z���������g�v0xY�X8
Z$X���t���Di�1�.�2�[ק�ݧlT��\���G;�s$ǋ�S	Q��2��H�	���Y΢e��}W=U�ߓĹ�	�oN4+��=Ĕ��}�Y��J�T궴%�3���x��t���]�27OQ�>�*�7�`0)ǽ���Jo:s���K��@��W�f�x��y�z90$�����ǿ�Ym�Z
e~�§�$�l$��\�
�lb�o-�l;w]>D�a&iMM��r�^�l^�	N���>.5�|H��o�.�� ѥ�}*����.������ɚ���-�o�]��&6�`�1��-��P]��k��.s�������P<�
���~��:O�6������.�<���?8�@W��@dg���n�F�{vl�b�d(�6l[�h}�8#�O@K��� e�'���$����-��M�(nv�b�"���R�[�~���gCSQ�Qsr��� QpL�S*H"�5�g�)����~����wlHO0�1�yZ��"F���@�'�o��9�]�o��Ij<�@?�Xyd�A�z�HF����C�����V�"�tч�ͬ���)s�n�g��6@9���}����1��	(�-] /�Nk
��߯n�?�!��8QL���\�dG��xx�z;��L{��aS$���|�2_֛޽��N_��/��5�o|=^7iz�8_1����f� w�#4��x39���z�)a�ڿ�$�t��wH��ƈ�7*�V�(�.Nn����Q���b[���ӿ�w"��.�vP�w���]���2� �v���\�V-*,e�=���]�s� ��8��;�#|�fߢ��t��;N[�C�ݐ�ܠ0?`�Ƌ0�wQ����"�M�<K~ޝ�}��"kn:�*-�'�����Z��5�����/���;�S��u�v\�my�!h���H�Ò?S��m��
1�����-%��v��>���0������q��֖0�Y�X.��f�{���N�%�@���"0n��_��$�V7�>��&����u3P�&�w9�I9�{�c\>�s��4O�·C��W��Fe�U!�V����Ȫ�av���GHN��T~�����g�����R��V��� ﯚN֝�v�7�</�=#�!$�[X���?�����ޘ�<`CJ��ú#�31Z�nD4�a���1�����*h�>^O��כ���K��^�V~�;�0�c 1`�w�Phi�%԰�V絹풦�����K��E�1�H�����W���nHJFUTk����0t}�Jn�EѸ�U��)�M4>�x@{` g4��%��xC����R��R��d!�t��c��d��["ᷱ�HK�޴ o�KM�uqK�� ������b��)�5��f{yK�b�K�g�j�����^��A�c��ȍ�C� H@���F���jѡ�VԀ��R���_����]�U�l��)��������dN�|���C�?�+G��9�W��61�jn�����V1�Z�G�ձ���hE	>C�ӫ�e2N���rw�o��s�RVQO���z�'w�]���Bk�{�?��=�Q=;����?��(Д7]n=H%�9ONϒ2��a�� �b� ��8Zi�p��^�v����#m�8�E.m)�Q�b2g��~S����>��evp�A_Z����r)Ó�?3z6�me���O��z��xn0|�*dE߇����0�r_��%�z<����#u!�~�;ۜ^�JF��X�"ҩ�v��ޣda��]��l����8t���F"�V�Zl�M;C&�9���{E���O��vjs����2L � ��7�v<��>��e��������9ݥ��+q&\�����V���7r�%�-�ѥ����ԉ��X�i���?Ü��.K�����J���ѯ\�Z4U���l�$P ֳ��O�O2�#�r9۬f�6��;>�xH=j�DR�)�h}MZ��C^�u�k�8��,l�����;Sߌ�����{�䟋EK�,�[	OSaGN_������TR�����S�@��6��Ow{��
��<�%c�<ޕ��|M;p#Ƥb���#�V� �,����+L�P嫯s��k��1a=,�JNcP>]��\'�.�A1J��u,���������/ˊ��q���o�.*/�co��[�Y�R��-�&�Vq�*h8�dcW����#Y��tX�ۂ�Jo�z��=�0�e
*&�S!�q�����$������k��4=|_��8T�c»����a䤒[W��Th=�}��;a�U$򡚘~N�HtRi�6m��ᬽ^c�z5g'?&f閑�OV���1�� 4mZ�+�2z%#B�BE���%��l���i��6�Iy�"�p!�W�b�J��Sܗ����ܶ6��݄f�i&��aõ��z_Hｰuzz'��k��6�9O�P�t��r%�Qd�|ƒAp����>�M���h��։B T�d�F���{|e�0f�$a��{�i)Rk��R�O�<wsYuC�IY�5P��34E�%X��#��9���^	�a
,s��b(�j%%�:��t���M�e���ݸ���qȕf�
�q�E�銘��~8���c#RcZ����QS1�YC�������W�8l҄gPxD����P2�6�+��voV)Wv�e��6a� �c���ܸ�b�]ƶ��U�þI,��>{{\ӟ�Ԯ¹��1)������oM�g��s�Jn�����^_mE���\L���D�G��s�wQz��8?:����`k��tu�8=!J�
��� b��3���KG��L	�8�z� �PK�t�lC>x�Ɛ�F^j������=�>d�z�B�S�0'�nm�2�+IU�a(�3�|��ͻ%֙�1qj�ƩW=Q�Zҋ%�A���:� p�]�;�v�}	�&��>���u��z��Ֆ{-���醦���Ax��U��_Ȅ\'�V��bu9�w	�Ab�u	�5�SzFT.�Ԅ~s5��l�O��o������,T%��$�Օķ���HA��;l�n����n�(hy3b��q��ﷻ�4���~G��2������ۑC��� �XR��	OC0�/nC$�I��^B��Bp���x1�JBe�So���Nqr 6��>!	O|�|�8����gN cy�<��D��J&�,B�D�iH9��3�%���G�61
'�e�T��
t[	S��D��=����8���N<f4���M�OFI5$mGx��{���R7�³k	�gϗ!W%��#��2C�0z�Zi�v�(y��z��/Wd%��@y��i°ȵ�ߔ��d�/:B0���e,$~�k��p�B�]����Q��Y�?����d����p h$���MSq�W�k�E�/`�;��TH쯂�N�����ǿ����S�Jp����+f=_����ݴ�Fzѝo�������:�)E��LN�&֌��{�n�1��M}����@��*1TƎ�,%���֍�]G?�|��1�p�z�9:��+J�b�Ӗ����G�Jv�f~�I����ټ$�v~ڿ,�"��mjs�����*_��N:��d�1�#?=|{�ڽu�9��e(��A�p����*�ۨ�����a�jv�Q;�.��7�B:�*h�mkO8�)�q��4�r�W����i8 @�	���\���{��yA��M˦�jDz�������1ʿq���=0�A�%%����BkU�����1�B@8z���@ԫQ?]MF��x���),x4�,+s��v�d}��G:�����@?�a/�~-W�OaW����s�����ϳ��$�:���o���h��9����g��&�Na����ho�� �ll�s���	�NO�p*mw�|Q|���`�� ���?z3+G5b�+6`W���y���
h>­N8>K�xJ�yQ`d��#<9�<��,��~��$/�f�b��Ts�P��^_�t�?��R�R�9�VB_�~?'G�(�s��X x��*�v�k�N�>$�[�pQ͚�D���ݪ�
�w�����܈	����품;��]h����N�2R��E^�������'�z�ffL�b��4�k��	�{}���G�rI���"O�lr��]�;��?8<;vߵ�
�Z{�og�˸G� Ѧ��V4���p�y�Ș��_���%����D��������{��2�5��{c=7��u��?9�F���J~8#�4TZ��z��)"x����_%!������aA�*��|"���
8"!��Jv�_�D��t��0���ņ�KК�1�֙z�A\�K�}�7�y��6����@Q�;T2�e��fM�	}7Y	U��UI���� *������BY��`,�L �ɇ&��i�}�e� ciu*!�\D�wԀP܀PT�6��1�'�5S!��x�,�gF"FiL���j<�|>��������N�q�-[^�&]&?R&�&R��N>ܐe܀�m�j~+�W��T�������+C�i3���;���>EقL�}K���p:��.
��K8g~���3�\=�����c��B}�$�5w3�9a���jOtc��p��P���
��s�p?�x�H��$t����k����TB�,��_2:��v�<נ�<��K�q3�見��2S�5H�����ʊzB�`M���v�F��z-�*����zl�u�=�HZM�Y�sc�����%�w]că�pb��D��s0D��`_�����{��W&X�y��n�
pdܑ�me���ٺ�R��Q󦉃��v�D2{xtq�u�L�I:�M�4�ޘ���A:�md=�s��s��Y�Y(nv*�<;��툚y�:T/U>ji����<�\��H>R`T3!��w�!�����d�Eb`dd��V���1f3����JJ������	���D6x����M�eVs''�b7�%��B]&铵$��6�ɓ���� :˺��V%=��)$8�5c��.:paϏ�6�K��:v�GgD��ms��;��|^����>õ^���6^����(�6�������=�������������j�g:�~ȊyDpkӃO�[�]�=X�r`�\��y["�m��zٞ�Y~�s�=�����-,AfTV��ʬx� ��V�5�����\�y~<�!$z)M$���w�hs?:J�h¶c��_LWߒk>�#���ri�<=/�:��OIM���T9O���׼�ZJa�NIH���o��r �}���xy�+�bEDDL�*ۣ�CC�cKɦB_�3�!��m�@6�n%��O*U��U^i)�e�������
�����w�.��HC�%�\�R��!�J]��XZjr*U��&���DK�k����^T'�ν��D.�k^�� �ũ����P�̭s����-��m'-�Eh��JE���B��㢊�G`��;gp������2H&0Pddd$O��\�`��g��[;=���a��]�X��B6f�ɕ�X9�,���B�e�R�]�.��������s�S}��h��#�C����འ�9�������n^^N�A��FT�k�?	���9|���Pbfw�p��4)x�����=��RP��(|Eظ�>%/kf����f,c��J�/����x�D�������l�#��2 ����=V����L�^����\�zNGG<�/�G<�xK9�ŏմ(�Ϣ��ClQ,���n���d.�`��ś�eai��Eް������s�3�=㯵b! �FU�Qn),@ӛ�\�sЍ�턌~�̑ܘ��SnC%���ŋ��j�v�:�`��$�U��-`hE`d<F}��X�y�hEc-hlą�8:9	ݼ��,=H%����z���|A�����!Q}�"A#$$��T{�l�a�jJj�F�`f�4i/$=��2�.P�Q!�e��E�z�No�Ҏ��Az@#Q��T��Ն��]`s+�8;-n�tum#$-^��m����>�ñ��.-�D�����	A}�HFs�!+�?P���K[�����򁶡���#s�1:X�����*���t�v��8[���!��3W����*^�k�V�h�:N�lw7u���oʎʞ5Y�ª;*��3E���- B���{�rmd���8����ZNl�t����;��Qҕ���d�B��$�b��!"� G���g�4~��2� �o�����\_qP_��[���^����HD0�U� P�1�>E����M�i�<�azT�����������Zo��:��;�!������e+	���[\��'[��R��ѱgg
���RRd�^�=�Dǔ۳S^��d��g̦�yV���������z�I*���8?F�)��c�Ϫ��� z�|߇���?�ump��8�r"!�p�ڊ&�Q!�wA]�{}�lm��:�6w���_Z�!��[>#��bʕ��c��Y��,.v[PQ �< | ����Bx��:_�Eb����S��B���l�jɭ���ҹE_����r3)�y�����]��N^�����ӈ��Ě�<%+��9���p>���������|��q��Mi,';щ������I^�'�^-'9"�	=JB�F�J#g(��d��Jr�mw�q~:�\��[�~u��Dӥ��y�0
R������Q�CsTf�^�(=+;��k^3�(�|5�S��,�^�Xx�};K�j�m]�mr���c5'�\m'A����P!����IE#��zv���=��[����$��������O.�^��Q$��J��^��	�_Z�>����U�)�(en̭��5��ڭE���4/9B���&X�˫�
qj9p���	xqo��At,���ˇ��:)=)��\:*�f�%9a��.֗<��rF��0��h_+J!;\��j!���1�t�����*!:A����!���h{z>���B���K쀱~2��c���wv���s���0^�%J��🜞^�_�u��U�hh���cH�~Wd���[I[Z�jؼ�������J��^��c��R~n\'$̯���!H�P��K]��C��'���Qo�ʁ�wfԬ�k����zRZ��9��_�?:"`�s���~�:GU �uѦ1�,_	H��j�,�����&��[��,�w:����aja��14�/��	�!���l_�^J��q�S�Ǐ���\E�#�F�-כT4ur��8�I��$W8�,�Ȟ��M��;ie��n&�6G��r��e/�/��:�t�T���Q5�5�P;4�sY��9��:��\��{|_s��~�5E��i�C%
�6vv�������R�T�MM��R\<<;p� Xؙ�ZYx�Ύ�ͨ��NB��n���&XBŝ��T*��ݢ�C��,U'��Tԅ�<�>��(t&����B�֢IJ8R4APY�� 6�����N���3�������"_M�-�v�1~�ų�B�{^5lҫUG���7}4�&e#�y�$�%�l�bC��A�I��6R�Oc�0Y1}�#�^�0��6����}>��|�   �YK+jaa!K�G9�i�����X��8O
?l������O����G=���|S����+�y�{��ḙ���T��O�[�kW�b7���<M������o��&��q tP����{4%`��s�W�"��Y��O�z�"�ݙB⿎γ]Z:c�o;�f]맏���!���޶���|�quh��z�[$x{�)��l�
ժ>]L�<��:x0����x����Ύ�[F_���,x�qp2�����Ip���W[~����[5�j�����J��YEv�a7���4%�R=n�F��s��/�#0�^9+[�ޔx����"TT[#�Wv��wGQ�E���K���k��ޱ�wV��.���c�z�~6b��΄体��Gk7��)(�Z!=���lͱU K.ujz:ddD������^�1�#<��-[E_LZN��'�D�n��:�_j	�!�Ǩ�w
����\-��ag����c��w�2��שIdX=��͐ֈ�N��x�T�q{[��u�V��mrPw�*Wj�6R���=F4m�7�q�W�G$�S�r#��Y�Ë��b�6������Ȃe�<>x���ł���'�j��e��ں�+�Z�0�͇H����36l�ʹP�K�����K�iψ�
L��'���ž��n+#�ϑ�%�_�t�3[�c]6~]�����|9�Z�	�+蹝�W�)�Ď��v��/����"���.���ໟ��L��p7IT����ʈ����%Ov��h9��x��p�K\�$8�É~(4��:aE�a�l\i����E���ՏO�;˫&��?1�� t��.f���@�vbUr�(��2)������k�1�c�������v>đj��J�y����]FfF��HxK���ܜ���t�:�P��w~�ӎ�T9F�n0�hUo�^N-I��i�x�b�D�`IO�3��) ^��Ak�x�d.�q5��nU�n�p�,'���H��{��Q���ߧ��1�I��Lnk'�\l,פ�0��q���7mH�|='��x~]�n��pt]A��\���3��m6����a2DvW�Y�dD��%���6����w���My_��6X؁�1����P�=����eh�O(	-�4�w"� p�|���.(��M�I9?r��"��EPG�@��I;�ů��� 87P���U�ڡ����=�c�6G�omaҾ^{]M��a��l+�¥�R-���[�$������nO;IC�7F�Z���]B����+���mwwww	��	�]�����ww�<@p��<�=|�����M�95̜3ջw����)������.�qs�I��\Ґ��w���"��h2�f��D�ӹ����=m.0�M��iæjQ�Y�G:)�q�FP�N3i{Y~S�6�z=�/�<�>_i��&2SA�{zu7�%�Z��]�05c��Wx������Q[˜�gFO.rp���r%lY���OG�ɏlg�{̗Ȱ�Q�}��I�0����|�+ɀ�_�̌�kt�"�Sh*�Bg�̣����2)*�F��L�  2�a�&�x���<�E��	����F
��z�Ϟ
O��<�J��9I�蚴l�@2��$�:���)4?tf�#s��rJ*nm�t_O�z�箿^]jhb�t��L�����~���u$�,�o���1���B������y�K��`u�������������s���jⲍ�����ݟ$eӅ*�Ë����-7|||1��6N��D���u��꺰�m=0��l��!�YOmS1�=��"�_r��p6��?�M�S37�������qހ��ɜKa)����Tbggګ2Ш�ÌW�X}�Abw��g"w�K���ۆ;d�E���o��x��e�M:%t��#�!����igm�����a��
�v���q�G��	r�|<[��lc�->I���C-55����8xF�+��?����Q#M��o��n�.v�5٣E}C8��U�T��8w�m��	2,:�[���}l~p�8z�P9��w(�yH;H`�DzTn���|�0����Bg��?Jb����e�˓X�y�`��85��_�p8l� w*��o�Ý�
'�}%]����I�f_L
� t�'��^J��s9��z�ږW����`�||�|�t�!�<�x���G�}z����Y����_?6'W��	�3z� ���%Y|� };,����Q��n�C߱k���Fc�*y����
ی�<7ڟ�����%>[�O�	��3�\�}�?o@�%$;��r3����>=�)[�}L��iZ�@�Sۆ"�#m�Rw�p���nIy����d�1w��
�t5�}�^��{�x������D@h�(f���;����%BNG���$P��h_�M��v~f�9j�y4�R���n�^�W����dK:|\�J��b)NZ��B�yM��v������2X��/�I,+_�i�n����E������6/��W�l�3����A[!��O)�v�h�s@��\a�>^�9/��(�e�H��u; ����|�5 Tq��E��B����
��J#��G
��z���ٟ�
��
�$O��F�-�*����MDjFw�Tm>�9���&>zƟH�0�w��$5��U�S%�C�� *���&��%�x�Vоb���T�X%W^�mj�k�cN����3W��2V�n�j�e����4�������(�Da�)��>�3�@A�s�^j�ұD��#�@���?���ٙ ���+��j.�L�/"��NcB���3���(b�:���.����Y-%̠rMmo�ꅂVߺ}ֆ�:�}��+��\5H:M�������=k�È���O�U�`��C��=� �Z�ky!��?	Ǩ?�[�����o>�;6겴�����:g�S���Q �� ��O����� ��ԸMm�/2����d�o�7�\��X�FI�.�b�Қ��5���&\�Cx������a��bC��L)��t�Z[I��|𶣕�\Ύ�P��iE>O]��!i�)��Ww��C��؉ �*F�h�?Z�]�ag'��m�V�#�3x�b��,E`歛<�(5���k@)�.�QqL�k_[��ɺ]�!>�)AV�X�k���r�HZEΎa$i|y�V�ى!�"Ob�V�>����mӣ
|�uj{A�Ϸ~"6���N-���m�c�G�����ⅹ9��B��r%z�D�����׏@y�K�(�;�5��Z����vϵ�`���r�AyU;~T!��`�ϑ\��!7���=�(Rk/T�%2�<lP}z�Ap�j��b�H����
��8��3��oM4�e̳�Ą�Uc��p�V������{�5����0�Nj��m9&.E�1��T��kyNk������'�z��#$�n��6�N����-�!F�󚠮iHV����e�,
���5un�y�L���cӝ����EJ�b����kZ<��w�"�˅��k�m]E�:�t�j���1ouF��A��r5MM8�?�$�LHX�5c"� ��M�&���X��Ҡ�|b��<��۟��fP�tx��S]���o���k}��Bh����'3�-������@+헝�e���M� �u%}������\���'c<���O.�x��!f���(�w�� u�}c��G27�IS��Uw��+��=t���A�,������	�W�����G�q�Ӌ�p�c�i0Q�O��]��о�T� ��md�\3���s����(�9m5��>IXd����Y���d�F����S.1o� $��|'�������w�Fi�H;�(��y�����%���������f���*��e&$���fވ�_�� x����Җ(��PNww��v]��s�\'777��,�zk) �	;��i�;�
��Ѡ�%N��J�}�v5�� �GRpxh���4���Y�H�]j����\vдXxt�h�Oe��Vs��q�?AN{k��iq�����+4nS��Y��ڶ�^��Rl�'�Dj
�8���?�X\I_>)����*}��K���}E�_;ֲݟ�N�|�u�w��v����i�Ae�n�,�_[�MY� ��*]���0����F�OvN�Xh͒"G�v#�z}�K����M}�x�:���:\�LޗF��g
��&�v��4ȣxq�p��s7���թ�����6��-�/^����o�d"H�}���0=/�ϊ�����[ ����o��?W$�/��O���qV�51�U��Cp[Gp�ى������A��=QB �غ��> B7����'�U�n=W����??�!�0)�ݸ5@�wY9!x�0l���1:H��l,�H��� �J�hn��~��������cn �O��M�4�3��5b��5�)2~,�	��`{�8��Jk"7��R:V;t�JW���B/�1?Km`Ѣ"�I���]��@R��g�S��۔����GE-�W�L4�z�%���z�����C$�Q��mthk�ed�[<�����4M:���H��7������(W�S������j��T%76J	:��"R��k3>}�e<u;�@C�eGG��3�;�ܖ��0����aa�Ez]A��ᛔܐ�r��%����TW�|
Re4�q���q@pl�e�͊Zs:ކ�u�!l� �N͎��FK�U�KIO�!���>�$R��gȺ�KL�tB��-+���^p-�&Rr��c����b
�[�X۶v?{���Ģ��,S��y�8)�u��	�v$�R�����<m�zs8QB��e�8�ę�p?hN���#!{�������&7%���zE,h�0�W��}�?�����.8��.�5h���3��C�C�ο�������z�ɩ"�k�f�2�!醾!=O���EШ�Q�Q���n?4�|�~գ����Y�r�C�~�]ÎF�{/�' ��.����-x��3���H1���}�_@��E���yqИ��+p�%��!ʏ�ի��}4��ݯ�W��>U ��)��v�o�z>c�U�W㑵��>]94�@��	�b�z���E���F��,��	�	�����I���T�8����`�?���/* �p�7B%�
D|t�&��In����ې��!r����{!!{�!x�4L�z��^�||��*�rz��E<ډ�7�Qz���.:
�<�ZZR"�����̃�O������ϳ�	絭nq֫?k՗>�c`<�M_K�^��'��vXwn_�d@�e筪��ϻ]���[m_ݞ���<�QH��9v�+�vW�����j�p�
@b߄|�A	��n�����f��2����@6����2)"ER�xe���;�j��s�|�Szs�C+��)��M���QZbk���(b&d�r��f�e|_������U4+x	�\X�W��X�"�.v�I��q٢����~�B./a�jp3M\���7�>�,4��teJ^�)��F~�7�5:)�4ut��D�#A��UU���F��!p�Yb����q-_�d^��
�	�p�T���sh?���`��tp1Po脚E���}�R6�SCL��1�J:Kt#O�~�[���E�ɠ�c5��2P����e������,�ාb߹�閭7sQ��!��Il�9b���A���*��GC$Ⲛ��� Bm���.H�P1RsZ0�b��o�J�@�)T{F��|��#��u�	ߣC��`�=�<��گ����6�򕶤D�^*�^y[|l��7>�͸���H���87�1�gd/����E�i�_6y����R�.��b���T�_Bp�4P�#Uf%$�r��aGbU�%!F�UoH�R����W�{K��8VX�VDL("Pn��ku�k�sǷ��Ya��m������BK|�Z���Y뱬(X���bnb�,�{Ǧ��ο�� �d�I)n°>�46�agt)��ށ�N�~�ƫr�Q/wJZ���}��W1�hѥ��EP�2kYfp�o�����^aQt�
<�U�	_�$%0�6�K��O|��Hγ��ư���n7X���I��Ƽ+�'	0�4~3��3K��j_�n2]�����e(��`"�s3�x��O��>�}���FU%�
¼�4�MT�e��䏇���q�9��*i���6����w�p�'3�Ψ1��N �P�g��lK}�F�����;  �K��	b��2���8D�c9��z�d<������?66v^{��U_�PbZ�v(^�*2e9#�h��Cgu=G�4:�x9�A�٧����ʋ�y�6�7Nz��B������q/
OF��>�B�%~�^��<�Y�=�|�~��E=9��r5.�@^Qu��{�Bmb�S{�/����O�&u��R�3s2�E���|k�sk\z޶g�Eav¤�����z[o��N�-�����Bo��y[f�N�L�/N�w�L�1}��;1l����r9�&u �Z������-�NN�C ��r�o�t�s��ح{�~`@�磫���:gKҿ�H�9۽=��i땧-��Ё��WZ?��j��9H�֬�������Y/M
�1>Np97a�^�IZ#�܂��)1��]߅\g<*�NF�i���ѥ���i���		��~2�D�)�|��O#�٥���g_p�!�{�?
xH�*mq���X	���ܯ��ٮ9$��f2vh<�B�x"o�&N�|����]H���Mτ"g�ھY��{t\�j��+݄���^۾{8lz�Ţ�����6���\ֈz��r`橰ߛ��a4���x3���w��f������|7��_x��Hm�Pj5LE�)3֣��bF��buQ���"��jI�t��a��jZ4$�_��L� �&��)@!��V���� jG���D��\W8�I�H�'O��J��P�k��Y��5&EJ5O}��XP>����4����GX�7�4�o3(=�<����&�ʽ��:�P�4/��`l�M�Ai����5��zϿB)�N�yWRKE�2��D���UA����!^�
��,�IL�U�L���AA�))>�:��O ͽj��������'EM��K��y\��z`i�]���jvB��I�H2���h)b���cU6�fI.:|���H�Qfǲ�ᗱ_P\`ɡ�q���J���%�#Ѻ��T�EZ38�����m���В�fu�4Y��;K��U�����<�A�V`5+�Z�Tq�g���-�0����|�3�%��sdddl�	�}��������2�H��� �/�DZ@�RH�_{j+84�vT'h�g�U�{�.��L���"|��O%b��R��x8$>�%��dUN���� _�y�4��i׉^����jk	K#���G���D����x�'����S�QP�G�zoTA>�S����W����Da�96>>�B�38c��J��P	
}��=9<
�P�E@΍�vƢ�w��	����D..[�T6��ZF��M�>Ԛ��30��/y���͸w����|�N�X�?��D���S�)���tݔT�t~�q�,P�_^M�d�q����p��Ɛ7�J�l�J�1�Fl΃���Q�Z�}sV��/��&���;�� ��V�C����A���֛LD�ԏZ^��`�v5�j�A��0��,���J=��>�I|^�]׿�49i #�yA��c�К�!���ԛ���mek29!��FWW��n-������d{�^C�
�M��d��d�L��C����]�[�3!@�������JPPP����D*����Y6�R�"�F-�O�p<�� ���ʽ�~������1��ߏ�@@A~��=�8��5��ɽH�w%�A���u�h�͝�s��8��Li+]گ��v\��Z:0���4t\9�e��y�;�!f"��n��Ҧ��M]co�΁�Qf�� IEe��^�%:���1���=v���P2�z���sR��,k�S���oi �7#�"5���yuS�����qk�h���l���b�2@Ĵ�/C=��͠�V�v%i�6�H�cه�Ͳ�� ��T|:I8��Ii�9�B^�ϲ W�����������#���1�s>����q�c���(�m�6��~����|�DlԈ��"��jw5f�ez/���;o�#K��ϊ�P��}<,''Ǆf��@�9���>8�6�儞�M�����9*﹗3�����������R��W��7�#���1���q`(�]��JB�_)�&�ƆtlJƒ�aLa�BC�\��$Zs#�s���9�ⵯ�3�Eޢq4Y�)�³6DTGe?`���p��ww+�����7Q�fЎ׻��1�9��%U%�1�ͰO����.$�Ќ�6n��~��37�9���t�w3�3�|���u�{��g���9�0����� ��i��>��i�D1DS�9n�!vc�:D|�gmm8���4�@�&Ad���dH��V���u�w�Avw�6���+	��*�Oϝv�ϞfV$�a�ӬT*;���w��3UD/0�Ư�
������-���a�������ׅ�i�O���g}B��G�DE�ϙ�t���u�)Ն���>���uKិ�	����ذ!�!���7�?M9��#����Ĭz��eк+���[��Zj�>f�\�9q>"�"|�`��UB��zOլ�#>�|�STDqh��������%��L
'ӛ�� /ݙQ`��������~?�*�Sd �]��KU�5�G���:�k�U�������?��!Z�a���Q��2/K�7����+(n��h!:�M��Ȱ�n����S:�_��Ϝ�'V������@����#�q��RQ���yО8�uC�NN�Di"O�K���O�:�q��ȟ��(����ơT���,����Դ�=]r�/(AHfFE<�����*3ȋ��t�<�la�;���XX��LL0x�������*���;!�}S�`v�@ Z v�U�q.����T?JL�]5|�d��c0,��PF��<#���� vX��w�\���=_�ؾ��ܒ5�ǳ;���v����"4��9@�	Qީ]��mJ_w��%�o�)�v���Dk� �DUB�	W����.ZY�0.������Ed����~ ����5Ʋ�e+�/V*�҅�>��2��Χ��v"u����8:x\����(@|u�����X��C:q����J;E�Ó�˱�]H��H�/��U�Ս<o�D���Y�t����t+��)Z{{;�W�do����ӞI2���7 ��כ���SnaM+h�wa{a��d+x`M�>M/��=`��|)�ʯ�1�%K����d�����g�b��ז
����]U�{PZ>?0-c|@.�M�%a\zVo���x�v��#��� �<�=�'�|�xUv����%�t)�[�Xֳ�~�'�I(����.h�64V+�XN�b̋zˈ�)���@!`��ŗA�x�:����`�;����贪���=�{���;vΒ�Z4�e���Lpp0drrr��<�N�{P ̎��zS�������Vq���PԿ�ݨ9B|���k��wg��3�TN�
z�-� ��7M[�+�����]��5f=60w�`�\6�B���K��y���	����w)%mIky���<j_ O��i�d�E��qU��@f��/��c��)����J����^$
���s��Zc����pq��Q��� �[�N�-|m
��x�$����<<vD_wE�nU�66��Ӕ($B��� #[)�뵬�VFCc��hZ��\��I�yV��>���b�Bs�ej����<9�P{|WP���B�͓�ǉq��9p9�5������\@O4��^�(�� <g k8�˧`�i���j'����)o?��(RM��f��$:����㛗��p�C�W]Ԯxk�G�n�����T���Zt�l���>�#]V_�hFae``>����kyz�{��v/���[��U��5���#�Ѣ�ȡwvv|�?](�����Ϳ���~gboo�ߛ�h���+_V^.�.b�����΋Ȅ)�0��|��X�~�p<-�Q���#پ�d�xr}E{P���H�ɱWH�6��Wi����'�$�Z�({#�/����!1�F���_���A�5��'>�!Htc'S�o�J8���H�)/���!�Tɸ	I���:�
z��ja��4����=};��aז�^~��V�ᗃ꒎�u�}���(L����Is4�D�&3\��%�����zZ���ӟ?�^�[���u��8�Pz�y<>2[4�8'd���c��`�a>]x{{{e��WG��!�9sF�}n�}ؕ1�Rh���BUW:"��X��A��d=�3k�� tLZ�${�8<�������F�E�)XhB&�'3�q��H�a�[�
M�k|y���54����z�������>�yv( %�؝cys���z�����C�����0N��sT��:���'��Y��*��GrYQ�_1��'Y���-h�R�����`���.j,$����I�U�lD/���M�!���L�'F��o��2B�u���T���j����5D�(ihH
HWNc��,�@�i=�tH�r'v�!�s�5�%�Y�f3Д���f��/>yj�&�8}���}��f���A�Ű�bئ蒨���K�sy�pB�3:���?�c�9]B�S ɝW6Dյ�:�G8��U�k��B#��>k`D������r't3x���c�������9��.�G~�Z͙����ɟ��^0��l��?B7\����/Y����s/�Ϋ���yd����:�.��10��Zn��ۓ8���F�3���|Dݟʍ�����S�u���p`;إzީV������	�Ԝ��w*�t��:*M�ƀ0�>��#�+��-@n�ED)�郵��v�9gU=ږD]y	�]Hl����g2�N��N,�QB���E��;�]��=���dȃ�,񙲑���Rj.PpF��5cr_N�����r|�����׶	�b�ֿ��٧��!/�^�Y��n���â>T�`pbbb�n>Eh����ˡ��(�O	�i�='�?Q`��D�2��ǑE��ڧT'7Pҫ&�h@�/0�PZk�<)�ӎ#7Ð��s�b�(���&"���� �6��'3�~_���U�,��h�f�!����8o��`!墁Y��H���X�Gd3o�eA�Tpq\���f=�j"�j	���4B�����{8nr1�4�.�����#��V<��s�9]����O_w�v�](�S�[���\����P�x��f��w�VW ���� Vw��}�^a����DJRF�n�*�0Bz'p���s��}�{#���)W���S���>p(�����;�k�%�<���q�œ�kz�!�^�8j��6L��*�����Q�W힮��<�R忷�K�Ka���^>����G4��lAϝ��FC�S�� MDFA�sh ��?�ぁc�l�����]g�$�����'���M���\�:� �1��������$��O/º׺�[H�]U��q�5�W��V�؋�,�tO9ִ�c28��m~2Q�"hHl���D��r��	/��Ps�[6E�c�����f�~��@�5i�u~{�7;���s�o�w�A���v�Ǎ��3n���Y7�>��MM�fQbCet���K�1EB ;��([}ٞQ��<��턉���)))��J�0�<۽��3�I~~yYs�.2��*f��_m);t�etl;D뉮�U�r�^�ȺsV׃�I�M{�`��0�k�t��ž7�'@�߯�ds�y�T$FR��*J¿�L$����E��%�B�N�1��_��?���=9������R�ԑ|�b������ѐ�D5��M��nGjU������������u��T1[B�eڟz�LDQ�ז��z��]ҡ�1�Ϋ�x�tʞ��_�����ڙ��]�v	�V�P|)N�H��<��p��#q|�d��2����t�gl}f*�j��X��������gE�%��Feuu�a�0q��W �aX��Qs�>c�f��p��:(7��-�w��59����JIO�a�"��^B����y55�>| ����S�?�ճ�V��Ċ�z�\��/�b�T?!�rN^E�H�Տ�a:I� �i�40�@~�Xŕ�d���Q�hs$�vb��Řl�e����)�w�y�Vg����K+�HZZ�K��j���3�X�SѨ���1��j<�(�u��2��� `������<����4�#FM��)h�T�x�g<�����!���)�F��!��z��Ly��QU%+M���,py�o��,3mS8��I��JU�?=�4	�8��"zLZB��W�:x�������q����^����i������)G����g�I�55!A�5�8�%S�+*T4���p�u
��-�UPPf�b��E�:<��(��jf�$�/���a��&�Kq3�����^��Z���6������� �u3�7���"����$lmTg{�OG���e��Z�y2�y�_��Q�q�qwx��$JB����n�+8�xՍb)�}�gT�F��k�>:w����Z���������w��ON�>�!�k����%�A4�=�����Ynn���~"df����(�#���؍Fa$o&V�3�	F�َ[��9���!:
��yo��y��0���|g�3���u�*�N�a��>Ƽ9/k����sS������3�ǁ�F���Q<h�.�=�nOX����y���;�'�{�	�u�]D�K�\$
�e�K��Z�*�z��j7! 5l�n2��ď��^;>�i���21_� �j�^ ��VS:7A^��r�3�7%�?}[�F8\Yʺ�TK��;f����a���%��5X�C)��{��_p���)�HG`��S�ۖ3�sE��[�䷴I��������Xtn���"�s<�҆��(��|=Q�!X�ń��q�l�����5C��tn�b,ŞE�=:�]��:2e�Qlh$�'?~^�-O�CeK}E9l�z2�~<�j�z#�jopF4fcbddd�^�J�_@>>���=*?Ñ��tzG�ab`�:;C�
$�2Q��4B??�o3��`�����4��E/8Y;ڠx~Qp�~{�#][�s��-v �Ƙ0F&��6;&k�b`L# �||�F���U�t#Q����ǧw��:{�y���-KjXtʂm�liv|�c�P��&��Ev��	��&N�ay�o8��*n`��.��#5ޠHxpn�I{���`L�Cx�����8��@�/v�Ah<��i
F��\�|,`��S~:l�T��%Pr�*&�:P�2����ôQ���j����[R�	$%���$͓+Nc\I_n��me���xC"��w��)����,���h�Ca����QW���8bU0jfY?�!:D��������=������9E:ં�H=5U�R3�>�����`�ʼ�N=�dO(ñ	��q �RkW9.�4]������r�����f�����e@W՚հ�i&�nEݣ����{��ڌ�2읙��������^v�)�9��n��y�h��Q_�-(��fT�5�Iho#0��x�'�n�إʦD��L�:�Xr��GHt��c�U����Z>V�~�ན�<�]E�K�r��pi����
e$�4đ^��K���js���>*�Wڕ�B���w�
��I8o��)0*���1�t�eX��2�$���/4�t)�K�_q߃5sJ>���.���������jXW�?�>�D�ؠ3t�(�"��uC,!r맰��
���UH��,F�g��\�R �Bk?}�ܓ����|�N�������_��T��o�5ۢ�(5�'"�t��U�[if�^B-|O��~�?�ǊzW��AtX�j��:��:��-������8��׵" j�(���Y?��鯇�,H�g��� -�����˞�j��Q�^M������P9����:��3��vG��
��*��r�ݦ�z�D��;V�.�ipl�R�zD��΅�7�tD�w!GH,p�eT��/v@}ϸ�O�nk�L�&��?�k�S?7�}<Ԩ�Y�XdN����l��-:�����<̾�"��G��%t�;r�̇�fp�V�oK*�b�;.�7��Rih�Ǧy*����_j-�U�@,��H5K4h�3&�!V����P�ˀ��^��"C�Jo6xć����y��Ҿ�~2mr��s�^��r?0OR�-�ܤ��;��9b���Ft�$�\��F��@L���J�M�JC?A��q/�7�7���6�ժ˥j�ء������*����M���	��_9-�P���-/j��v��Ư�����Z���<s�kD(�@��p�:}�5�sE5���\"z�V�B��éu~�Y1dTIj���Nv�v}�f�</�nO'8H��.�g�}�S�6_�L�Q�I���c��O��;��=�:k��Hd���x�yu7��;LKe���@�TӍ�۲2�`�4AZ����~�,�;=��Ǹ�����%�	�x:BZ[�.�Yp�Y�#c'[�L�/AJ��H�g!%{�޴���x���	�ZF��������ŧ�2~	|ݗ;�Wq���'����&���)�=��&숃˺���r�������kד�����N�;�<�]&]��kؕ�������j0Mf�Ө����o�+��_7"�6ɪ��>PxN)����z���=�W�r��<�:�:�N,-��l�V����.a����ŇCR֭]�Z�v+�2P<�SGYƕT�����d	�#�;<s��nu��/��(i,TA��P_	��y�jV�`9(�9w�|nC��7�깂:<�y�����F_zot����(�s�a�4iJ9�{�C���fe����G���;��W �=s��o��pD��{q7��oGz��>\Xv�zY���i6#��6�}M��7C=�X�z�i�}	�L��C�,�.R�@��I�"~Ґٰ�s��mU����:zh�������Y�Ы�Ԟa��fD��$��r����}�*�~SQ�Ϊ#� ����9�(w��GU�F�L���9��'N�f������߽�����[�ڝ5�CPX;`N5�b�㢻u�ek� �*��;��%�����j+��z�k  �����/M�a6���U84.��g��/�{=�	|�6yF#w��2z\�ş~�T��R'��I���Pz"�AH$�1�H��/�8,ںF( �����E�O�)�^�6�U�	�;��k(_�M�3$J|e���d�[NVd�-|]k����u5Q����s�)���P��;uD��Uj��5��v?���n����ا��[�RS�7|A	��1k{Cd�ޓD���s*4L|خ��q�؍2�cC�V�y:��6��+����k>�b�G��)�hh$(��WC/�����Y{�,���)ښ�q��t@Xkf:�i�P]{��o{�*:�|@�?��>��:h�*�v��l�h����cGZ��տ 3�'�,���F�Q�ۼ�����x^�p���nE�8���c�`m���Y������X��C{�ř����[�&��T�����틳X#�O"��%3��+*X�㵩�ڿoۏ~����5b�`D�U�������<:���[�x�^�{R��.�����ѹ; p�o��5�����WO�����Yv1f�_��,Hx���V�f��������x�tL���2-lX>x�W\�^�M$\1���>&��J�L_l��&�f�'1$������=�P��0��~)]a$.c}(����ȻmV.o������v��#J�!����:��M�o�o���||	f5n�B7%����i��}Y������iv�MD�7�O�V,�Q�4��mڢ���@6��wֈ$D��&Sjm���1������`9�S��l���1�g�'���4�$� ���wK�y[C�~�o�`[دܱ�~�?��D��y���j*vԜ�e�t��8'��s���J5~��޲=v\���~uI�K֊�O]@����u���G��$;�x���_�!Z{B|�������TPK�$����΃�y��d�i�:��R�O�xlwzL��S���~b8��]5���2P5��b|���Y��lX�ST_K>A�Ɂ�+�
]��f�
��FdK`u��|
f��hg�B����l���E^_7�[�\��xz�H���:���^j4��k���s�g~f`N��Z�^���´��r�G��JU뾢��D:S��;{�4�]�B� �3���p�[Y��&�j۔Q����O�VyT�yt�e�x�x�jl�3F��{������ߥ�s5ǟs��	���P{�ޢE�c��9Mf��z����f���/�[+p��A��Szaw?��A�pa���n�ƶ>���i�V\����o'�k�E�W�&��e����)N(�d�Q�rL�Gk_5s�iI�=}�載`�`�E,�N�%��]tw��矶��Z��_&8���<g��[^@5�I���O~�t�6O��찶�\��=}���7����uq��o߷t�B5�z% 8?_Rk�}��)�c�ZG�1�����`=̇G�\�=6-����"�?���[��ݗ�h'�/�M�_B�h�N_�����A���Uu�T����"
y[Ջv�iI�w�b��g�堙���g>Oo��kM>ʇ(t�����t9^�"�k�52�o�y��?`
�?�q��K�)��S������.&<��0]�KB��L�Q�ve�Y�����ԸC(5�g��Y-fTpN�@79������xg؉��%V������6�=���h)XǢ�=��*P�}�ir}�$b� ��e�\�3a�ץoG�/�R���/�'=����9��ɓ1l��N�X���7SO]��j�p�6�j%����2�T��W�?��G����I������bF�nzH�';�!Lh�i��:m{�D��M�,my=!*y��x"�v�/�:T���,�;����4���YҞ���p6�mo���o�z��[+��˱�&n^����M;���/$0��B�b�C'[}�.��Q�2���πS��j#oB8���N��~�S�p��xǒ"K�p�M����XjD�����6̑[{�Q,����M�����<3�\���@|����������N��*\�(������R��gC(�J�3�d9�T�~�U2�l��/D�?�5w �GS��{x���69��۲Vdol��d�qS��P��RCX����HW�o8�7�=*	����W�>���b$*wpr�}_u���QE2-�Y�z*f���8V�Q�&�f?���OǗ���d��4�Dsz�%Ζ}�Af�_/�#�S����R=���+���F&��1fx�YДe��tF�FĂ�/����:�ܤ�@=υh�FF��=μ��6O�r��}�Z<D8�S���5'Th�3-��	�tǾ@�d����LpWD��ՙ	��)k�H1�	m{��cWr�u_{���N<��+6�l��xw�[g%Y�k.�VR��V��&|�<d�Ώ�U������D-*1�<�,#�7�t4�y0�a���ʲN|u�lI5��lL��~����ͭO]	���S��>��V��=E��m�Z��}68Ǭ6L�}�����a-_$F�3��W�Z�g� ����+-�T�$R&xH~_�$�@h�!iQ�e�Z6v3GJ'좊���WҢ��m���{����-ܠ����{�*��Yˮ�:�)����Ӊ�?��K���芡��ۭ�,����� zy.�@� ��Gs�+C�b����[�hf�x=qZ��^]�'�/�$����}Z�_b=
�I�ژ,}{>`���TT�cnКɃʿ�|n������L�R'�P{��o�]_+Z�AQ��7�ny��s���t�Ã;���!�wwwww����݃�&�������'�+����a�T�޽W����>5��b7���Z?g�켯>m}�$;l��G��qo�O4;�E#>��r[>��w_�h��b"�Q�C [��[ٻQ�D��⯖W%��u�n�h��	�O���G���D�Y��R{ �,~p��۲���z�Ğ�W,]��=w}����{�f�W�]Ix��6���U[��5���gN�!6=���D���\��� ��O�I�@ű6y #��n������60P>�wt�F	�!�j裂(�P��;�D���ި�������\Kџn��,��u.]�q�f=���=7�fQ8@D��A#������t�}rq�U"�	��1�/��a7����l'�3�_�ZGn{y؟?H�}o���u���@�/B$<�r�m$��½���Ih%ڳq����%�ɢK�43�m�y ��+����m�v�/��X�Kc LS�=���hIG>Ǹ �j���>�Vs�����-[�SJ}4f���w��ݬ�00�&����ȑcH8}���B���&M�����&D�9q� �~�Ȣo*j�Y��df׷�K������zv�:��]יh��!�z%���)��v������p4��<.��YD@E�(}j��y�ג3��s� ��d0]�q��BF�tq�XSe�s���1a��J~c�'�]l}�=�jh�(�n��j� ��c ����$���,Z> r�Y����m�?�l��3���$ad�;�aQ�w *�e�>��Z�� ��~R���1|dr�}�)onx�?��^��Ȼ�T}߽��+]���'Տ۱�b��s����!���m��(���pZ�u�e�H�9�W[�F�P�������JB���N�3����7"�I��6Cn4y��n�G�8�|�y��|q�a�.�y˸'^��Ԏ��{��о�VB�M�hb�`��}2�6SU�u�1 l4��h��%�{�>���2m�Hc�l��F����F9+���̲����d 	~�̫�3�"ȝ08/�Z	���ʱ��W�OZ!.W������W�Y��I�f���H���@A��T��#iz�k�t$�����eVPh�y��\ �%l��h$����?V����	�j�B%4���z>�U2�M��9��XI��i��m\�x�:����Ā0��m�hv����⺦��O� �]&��~=Y��f7��X,�:s(��&�i���؜��#��:��"�*ǫ�OK�>�O�͸����ZI���>J�݂@5�x�6��J�^J�\�K"�1�e�M�
c0_�j3�^����V_�D�	S�7J�1R��ń�]&D�q��ڥ��jrw,��t��|�r�������sPҎ,(�u&�	�c�DM�j{Q`���wt��a]i����j��[Eؕ��+QVÎ�Lr$U�~Qm$΁�V��U %"3#��o��Q$.�Ly��bƠ$@��2��l(!��a���;�c;fN���}��'��LN�ciwÁ�������@G��~�jO�7ƚʬ��P�>.�_�r�j؈yz5,�͟Vw����$�{�T����Yߖ���,#"�l��m��2��o!.�ӌ��G��,rOW�2+�P���jԦ#�V:��j�zЮ�R��}��&�(k���k���\�s����5��'_i��Y7�mI�R\/9�F��>V���>�P̿����x5��	0�	(�{w�$	��Go=��*O�y��>j$	`9�"M��̼p��D�ˋ Q�Or��QR&���3�â~�p�d�V� 0:�Bo�[�h
>4{$@'�F����|:�>:V8K��{n�׆:g>qz�By`�>�^a٧+�q]����[�G�GM�IR}��G]8Tl�����ߤh(�Q���U�"a�1�F���PB�p�e:+q�j؅J�����Ћ++G�
Nf�Y�5*�3<&��p_tɍ���U�*��mMvS��k�>��I��u}p�
n�Vt���Aa���]&Lц�GC�:%d�Y��;��˷�������{w�z�
��O\ywJ�o��3f�������#���#���pj�Kt>��f��\�P�X�L���zҥj���YY��1�,��L�4f�cG�͞��!�7#�m���& �`?)�!ڜ�1?v[�,�Y�Z�
�<�ƴ�y�:t�7��/8k���M���p���**(��CF/�q}���O�)ID�M/���Ǜs��A�&���Jo#$�]��($	��ݻY9��$���n դ�IE�sC�O��q��q糶�49������� ���9�?0���x���������z�N� C�Y�p�����I��~{wYY���r̰qд�-�K���F�ۥ����ok�߸�n���ͬE��k� b܇�%!��OIR�ifb�]� M��F��c�
�T�fs�$@�iXM��7T<>Hy�2�d"B�.T�~���;�:[:�������3��$���H�Vpp�]H���=%wOFR 0ٰ�
�u�yv7��j�#J��Ng��I�st�륈De��ԝ�L��X$5���������� 9 \�X�
�Y��0���})�++D��/l��֪&̡L�Ύ����7� �cD	;m�ޖ	w]��)��%׍b׹ݣׇk��
�\��e�� �@�Rw#33Jq��Y6vv��Y.;Εxq
J�Z@A�p>�|��g��"C
���#@�<<��-2@�k��y��{�NdEx������=2[��>�"���U���\�;g=��^9p�.Vn^v|��U�*��v̅��SU�)E�$.j��g,Dl_�|������(Oxb?fL/�s.�����jI��=�����S����9v��1�~C I��uWǷ�g�ӎxZ�����fe %�����`Aj�s@��8���&��#�ƪ�pnC���tQۀ@b@�'hȓz����_�Rc�����\��6��~�C��6�7jY����\�0Km��^���o�FG�'@`��~E>2�U������n����?�;�f%,l���OU����_����T��~2����'�AG���Kf+ʣ�ҋ܆�cS�����I��%����j�f���������1]4d�N��+q
����&n0�ҙϹ|sӃ�̹�tQ��V��W��>6\���zCy7?2�rn V��?B�ў���aь��E&͗q��]ӫ:�@��5?	�I�L���>r���\se����q����@E(�`Xf�J" yQ��j $u�}_�t����QϏ���ŝ*}X�H��e������&z�eii|2ev+`zj�ב6���j�+�έ��vB�iw�&��s�ᣀ�H����'�q��Y�A��}�YXu�Q�v�;A�x�Y�����1�f�+\ ���	;,ܞ#��+�˶�}����6�
1�t��Z����M%�d�ڷ1:���2�2�X�W�#k �UO�rjk�*.�fJO�
Ñ7W"� ]�0�k-�= P�?� � �O�=��O���cwY��6��̗���R��V�Kx�h�[=5�Ѽ ���>�d_�+�Y����Mӄ~sC����<�:MیnÅ�$��';U�����y#6$]t�8��4kP�R-j��g����PWCS�����;�����l�<V��vsJ���b�G�)��h
?����MU�)r��P~92(7��xbOԓ�7���(0��2H�|$�Җ�i~�����^!e����	566����O�~fH)P��O������V��6�����@�f����Q]�ME�ܑ��η��L�A�<�Rp�Rm�Q�@�
LQW=I�T��|��y�n�����yk)v�i.&�s 󱷋���:�������tA3��8�>!*�Ĩf��p[�J��N�Ξ�͞6���t�3e��#ƚ�T�I��m�ًf�v~��C���w=���Ҧ��ug�C-)݄Hv?SN:_�-�s�Ud����~O��ܞPp��z]�(v��Ŗ��ǳ�s*��<��5����4iVm�5���'�����C@t�JA�Ƿ�-����NK�7׭���Y���eS,�@����}��$3@�p�_Y�>����5�����5ɢ)L��\�d��3ڣ��� ��ᷴ;���0 r���,te�N�8�}?���5�0�5�2��} �=J��y=�y�b��vM놻ǡ*e��#����M���J�40�	�9�4�žzt�A(��!���={t'�qfw��{��M�
�-��_m#D<?�1��MpTE��44�~�`�R^p��I�w�\dB~ȝ=�Wý^���c���!��+�VQ&���bv�1�����#b�,^����t?�ǆ�&�a���K�WE&&h�l5����U  ���q 9U_�M�`
�ؚӑ��'�]L�'aU��f��\�����*�'�2\`^`$�w��>:E4u:��-�L$�F�--S�6���z��~���!�A��=����)xʴn�ɕz�����0P��I��~��˥\�n�K�4���`� ��k��e"z���{���'��͆zW�A�]�N��U%�O�2�Z�Q��(b8���In17{�1�G���_ T�yB�8o�L��s�g�!m�B�����Hq�E�T�_Ru��t{!o^����ե�G)Ä����BA]+A�Ct�M2pE#FX����(~�˴���s�bQ�-���׀� �
�����?280[;�c�G������
�h(��p��D�o��2���U��T���T��)�e�P��\iݹ�S�`����QN�"�Ӕ� y�ڇq��җ��ZDT� �'���őۏ'��� �'�L��^XȄ��cFQJ���5s����R=����	-��~@]56��.���bd&��(fE���Y�@��F�@ ���UƯ�#�.j@��
&4���w�߽c;��˓��'-c�w�a`BDb,:a�?�3���y�W������+�*�'EJA�6dEQVW�a�Y�(�aN��j��*�~d2�t�h�R*ּFV�W~q~�HOvx�I7��'v��i�0I��`�U��A��7ɿKY ��q��~'2E ���;�EM{3��������&{�.sƮ�e(��@xT��@�C������;��4���SI%WP���F]zZ�5L�_k+z��N%~�3A��[�8�{M܂�x�k �¯2RpJ���X}���XW�d���e|+�W�����_w�I���/�=B����˩�C�\�*���ږ���by3�œz 1l�@�4�@%2Z�a{�|�gU�}]�ݷ��$D�2DD�;,�D&E%�^m��wD:��u��m�����&U� �'K7�����23�z}5�h�(���^)]��[��'`����{����m����9a�j�՞�����/���/��u��-ϖ�lQ`��|���8��9�x��BL�P�4�.�x� ކQF�JN�5�U�<%죙U����]�"�� iN��C�5�n�u,ځ����.eD�˩���y�F[����OV���TM˄ԎO��]�7{k��T������Z��I�4{�!]�7�k[s�M��0Nd��/|>�k�G��1Fs�Q{�&\	'�
����T���&�_����:y���:�9���n[��t���5J��a��dS�XǼzA��{��Q���!!_��?����U/�����!���ҵ�U��Ϯ�LmQ�ĝ港�/�T�ZoX3�h���M�
�(��V5g*�iw+��Ř$G����P��F���`t>�`��;����A�奄�����t�x5</Κ��KX�z���F;|9+���*���f��	k�e��W�2�Y�ʺ>�Q��x��.+ף�)
D���Sz�����fP]�=O���ּ�;��1-�;^/t����W��<�w�=`"J�4��r������!BMA��B���������J�$w�	�?�iW|��a�kj�x�j�EX����9>�������7�i^G3��i]�0Epeg�q��V���p���փ��%/�:[eg�<��;�o�7�1�E����_e1n/��5S�V���*1���ԛJϹSB_<喚2�S�"��>�!؂8�9U:Ci(~DEZ��V���k����W�,q�R$��u����62t?����Y,�����]ɐ�e��u1UW0�m4�QR��������k満�/R���	�}H�H�������߀�i��Q�d�0��F�"
�L��a'b1 ߸�|�C�I76Ҳ��N\\շh 0����qft��O�~�VOar��Qj((xtt�Y�=���H�Ï(���0Y�D##�9?:��!�w��������kr�Y��
�������HD����u���p������~XcM��ˆ�]Ƣ��5��k����v"��5uT{��Q��_4č��:CŁ�I^\3��b�UA\�W���0f_M>y�_�c���?�~�byRc���Z���_�m0 ��c�hR�~f-w_[���m�βC ���f����w��z����Dx�4��9�¾j�,�h���a��`���pH(��"8i��A"ZW�*��&7��|��Q�D����L�23o�D��M��D=�xFˎ`��N��Hw��8��<�B*�olɔ�PT�l��Zs/�0�-�-�}�+6�-17�ˁ� O5	H1��B޸�!Vm�+�]B_Íᱟ[����o�Y�5��o<@�X��}@s?r�ˢZ[3L�#y�hzV6��.�`�c�NY�#)Vp?y�豂΍L�K��8%:��S�\H�l^IЖ�(��Iu�6�f����5�`d�JY=��P?-��Y�ym\��R���+\�O|����x�x���"����p������o3la"P�����/TQƽHIΣd�W�ح�Ș�1U���Cd�e��� ���`�.x�B�U_�b�9��Z{����y��z�z�.�d����Y��@�?G
���u|�VO�CUGЦ$�*Y���}{m�����[�ǂ�;�5$Hm��ڢ d�}�>D1�,`6���3� ��(? ,�h�hvˢ���F�e]�aH�\�������|�,���
maaS��<y�IU.��������0v5_���ݧ�d	q�9v$R|drqӒ�x:A�� Y���1��(u�R���.S�:��Ҿ���4W�Y���Cl�EVF
�U��^�,;�a�����"e���~r�D�X�E�0x��1Fb��xvA�	�֭�&�R�Cʫ�I��ԏ��C���h(J�<4?�O���,�t�90	�,�3n�SVY	�f�����v� ��͏+)��DB��:�0x�s����хQ1t+�V�YVl.�4fO������RQe/�w@��2��@�ؠg���s�s��|Q��y�PɊ�w^9:�ve��´�2z��2����y�߁���9l�0�K؞��
˜�,���ۈRW6���:R!Rd�qqj��IX1x�ߧL��PN8#o��AV3����4#+}��`�iW������ks��z��L�f��PR�A�6���a��zl�1iۡ�[9NଔQ�?�
6�0cL���y+��I�jd<=xTgt�	�XS)�����nI�Ľͻ���(�P�X��DF&�?���b&A\=���S����}��4��s6ZA@Cq�����S��~�ȧ����}�y匑�"K���䁫�P�Y+�%y��gsU�,y��'W���	^���+]�A�s+�(;@h[��5�]��-����[.����
����t5��a(CL�^'��	kL-�u��$h��#��j��g���:{�p��h��?�ׅ��P����kIL#M1�Ч���g��[MG�f�:���3�����]���6�<��E2
v�R@�;�N�4��~�WM9��PK�qG$�u���0@�`3Y.%7����zt�yd���-'n����4bO��A�Gԝ���*pG]�tD�a
P8:�@����ɤ�mg��@)U��	�^�ՉJ.җb3ԟp���5����[q�6G.�6�&����ܔ���Mn��������M�dV�y/�E�b�/t9�$W��Fz� �+�=�I��v����H/����94�TC�}���i������{��G���6�{`�|��W�	헠����!/"i�c�>�*Z*�w�%Vk�
q���d�L��{p�n��`Q�C���4��dɠ�Q#�{�s]0YA�7�)!na���«>r��bG�KX�.E�~�1�+ �O����͟j��=&�j�9W��D�|7��Ф(�����s/t�
NA�9�S���)��>�[�lu��o���ڍ�bo�wV�?o�/�{�U�����z�.��>̮{���5E��n���"7Ҧ��r�#�#Kj���韖���P��u�˥�H�v/_���uh����m���t�`hP)�#�]4�z����{<�����8���V�}�����p��4��c)5���HfQ+r(!�J��</��O��?��_��;��
퐌��w��J����i��.��H�X.z�<���U͆���y�����6	��m�K��.��NGc�%=��u������ �t�%7A��ZÍ{6�Q
z6N�`����@�J �E}�L���jӛ���,�㬛if�I�T��Z]tb���v���×��ڶM��9����=��{2$�����
)��|L	�_x�8�ѷ[9k���Ev�M2�h
��-�5����Z��KpyE���t��C�c]��}��� �A��/�>\�����C*S�ʯ����)�;p�~m�A8u桝�6£��W�Ȳ������T�t);z�,+��O���������SC���iנ��JE�l�Q��9޶8��{�wͯ~]tf[�e���f	1�^�)�z��'�Vm�
=@^��g�P��6���^��c�:v���kt�~$7�(yE!�$�4& ������K��(����ӳ1wo�C�}�j�'����!F��6s'/���FًJ����_��	��#���7�E| p���kpr�ә�!<��I�������8��R�v�b/��N��p��	g��9ݔ��BW��B�-��jQUɡ^K���ij��#��ֳ�掠�i�P'��?MmE�ɬz.H���{
&M!V�Ԁ�
�ޤJ1�Ox��y]윪��o܃*�q~hu���G���h�_��s2��I(G�~]p���l95g�ѷ~�f�Ao���d�}�����t��Ty�d=i'��
D�����~�Ot���m�5�3C�0~�Ӡ	����E_��q���������J(@X���C��Q��������э�RL�{�pR�?�m����z�	F�l�<g��Y�:b��z�,��z��ϟIٻ����W�l
RfC'N��n��l�O�|q=���9�'�_(���x�E�^��=�}����)M�&�>��V����pc�}$����]�,k�O�f	��PHEz^��k�%|*����	ȗ>=:��4y��9m3$��+P�tH��0��F73ڕvB��r�nZ�Z�?A�R�۞��~-ׇ�����hQ���/D���F������c �4����A���a��*"m����,���r��3~K��t��IZ�.�^�5�d�r�y�U<�cx�-!�����³���/��ll���[�;ރ+�����/���h������/��+S��u��8���|��vNS�����e�K\	^��]Dq+�m�A-�3�1�8��H�hd�����'�cRIW��w��&�������Kb?�^M�5mO_�?Ś��'������I۪�������<��惋�J�
����^�J�q�[�Ŵr��B��[al�r��Wv���ۧ(sי)��?~��M�#�U��ik�*W��_^+U� b�F�#`�n�s,Oy�ӽ�����r�K�"ZAʼ��9(z��� �!}TQһ�K��n��E��e�@�y:W�������~��{v����n�����Xyϻ�3�� f�.�um'��ٿw�����7���Q���UZ��߰�������b���c�#qt�
�~�&�u�&�4b%���u}ǣ��:��s4���Q���ٮ� �1y�+�s���[�<��Y�Y)�Zc����*�᠙��� �:z��N�;��Ңc��ID��Ƿ��7Iy܎h�7�~�7GT�B�q��D����z|)��<_��O~{|٘�!e޽��KB��9�*�_�'���.�|�d�NԺe��0Ns51���S׹���ϫar��
�T��h
��h�l�i���y��4q�8w
^6��o+#����w����V}Z�	k���v���Z4m#���+=e�������̪#�#���/��|}ص�4�x<�G��
T$|f�s�z�2M	���t�����%�����Qҧ�A���MQmJ֣E~jаF,�;��nq?H��K�f��#k���.��E�G�p��ǿS̢�}��4�=�%��9�'�sEm7&�n�MP)���M�nF��p )/�(~h�k��*����FP�-h��B^D�!��ɧ�k���� e���l�A٩�7B���a�N��_�Ub�f��l� ��Oo�\��v>*��h��.��>?"�܄�b��y[�p�����Q|�(_��7����3�=�?�iy��zo`�i�Ik��:1��h���Db��G���8�_��nΐ%���q���������p����:� S����L�ó��$�?����hkϻ�x�󬭷KG /���U�M�L��q�8j��EHv������k%��X�>N��@[L�fRB�J�K"8��qM�*Mx�����mܫ1i�a#�i���[T҃��;z�o��j!)K���1��f��;���U��t�>	�Ed!�i�U�����VR���aV�$2�@8��+}#]u�-]n�����Y��!O�G�)o�����v���p���&o��[�a?ҭ�q�1����9���N�5ѵ��C��6�Y>`��~-�[Qn En�O�[&��I�!���*���&f��?k";��Os�Wr�x�/���DL��7uC�!�2�yLa���pNU���E0ϛ��T�޿�*��>��-x�`\�}������qN�x��	,��ߧ=	�L�E��u�p��-^t�Mw��f����ز�]���_G����"�E�C�Δ��7Oã��+�J��?�[�K�Y�4���xp��ٗ��[a���R#��xB�/R����I�/���L�Oa���&~ ��j Y��C_�HH��N����2b�$�oV �*3��s`�Ê�C�UW�7,�x�=��!���?���jzlx��L*ZK
�+��bv.GZ�-F��Qg�e	�oƧ+��+[b#�(�C}H���6K�)*'�gb4���CA��q�\%Pj��TE�ol�����D��(�����h������i��� �m����14QV��Ens�����à�v|ﮠ�����G1�����+�������}u5��K���ٛ��n�����&�ؓ�odu�&��2�H��%��� �!�p�.:kѰ�ܨY%�u{�3��̰e1Itl��3��k?��MTa0���. Z�n����U���p�T�=����W
Z>
�	�#�o����;-8��=��&D�(O����V�� ���ϡ��E�I$��1���CEIt�z� a�r���H�F��5br��.����Q?���
�Ec��:�<�"R�zC5Um�p�Cd-��o
��7;��k9~����6�����փ�]��r�C�`\ �'����`t%ߟXV�kUU'^-u�ΝOi�n��Yx����\DT
�dn�U�,�X��]s�FN��$��!`�;�q-➛s����_�w���mMF��տ~R�ߠ �ˊi,$��U�N����K��B�c>]  �V��E�E#�l����_��i�&�΅�8�!06��Qt������>����M��C9-�ZY2����6]��m �*������bh����,��>'�Oz���z�$�'�"��ʣͰ�:�T�r	%8�Z���ZS�W9t}��LU�k>[s��{���|Sl?7���6�xH���cS�/���6�!����<�@����©z4.�K�����"/M�.Eᵪ����L�f�V��1����$t���rr���s���1y��'�dG�Wܿ�3�ض��b�A�jn�Y
kZ�df��p�5�6���;�fɋ�>��u�x3!��d7���)uրן�kg*�����(贵�v_�p�`�s/mg�z/�WUG�[�h4�MPh�D܀�{P�7!_��O��^�?O�W'ְD�wa��u���rvy(���y���HpbV4����ן&?G߬�a�@�&e�`�W�IG�1�u)��1��,�S
�^��`+^��%i�St�<ɸ`Pe\��|Q��7p��d hj�wi?��i��@(���y�0����g�x�5�\��V12�_�Fl,svw���D�_	�s�T�"�����7%�T�VS��v�U1�e���ϝ�Z��5+�Q�01����Z�8�H��BV�I��^��M��?�K�;��Nψ� �y���6�F����p��ʜ��-�\�
R�_��b��aퟣE��d%����q0H,~�p��K,���h�ݠ�(��A�o:N\`�8��W�Z��~����՝}�yk���(a	���@�_�7�	��g;���L՜�5es����E�6?��$S��`TwIS����GW<ϗR}ő ��L&��Y�T��4���Px}�� ��,�t�����#�o!ms``����հ�Ͳ���p�u��w�2��E��I��JL�Y��g�k����K8&����H� � ok/��,X�d���M:�(|�b׏z-�WЉ�Z;��!��T��p�DqHh���Y~c��>�r�<y��r���=�}�b?�qd�YJ�n�i�x4����U�6+T�B����_�6���/����r�#�Ut#>mWOӹg7☨6�=���"���3 ĕ����s�c�}I�N�PǞ�}��Gz�� w��1�r���H+�<�,�����kP%T|��g� ��}���bfj�{�D�$}�>�7?��=V�b:�g[�h���Y*�)@�=�exr*�څx0N�7t�j:��VH�; �│���m[�_xx��sN3b�t���$�K�Y��D���p�E[�G;zJ��@��ӌ��mZF�-�/�g�X�M��Dԯ߶���z�7?;j���N��}��as��p�^>,a8�-MX�ڲQ�,��S�:�O.U�<��p���̔\!p�C���wZg����AQ�n���Ǣ��."@��o�]�t)*�p�]ғe�.-i��?%�m����5`�!��i�F2xv{��%	��M���Aū�����3q*��e�|cl1��\��]��I�x��y�w��K��H��9�m���1�r�B��:���p!b�}-�"~b3e�����C C_
�g��/�~�i���$B�1� �M<}IsP5 � cb��7V8���׸~��g?<��^A���V�/B*��V��}�q�MyIc0À�<UD56��/-ͻF�y<��n ��HI���֙��o��z4�ᵢ�y�����)��O�p��������ǜ�����9bb�7�2���׮��!��v��J���5`�$�m��L��H��������������,Hxri�u}f1��Y����0v��z������J��9����)�%t��;�J�=w�&*�G�&���9�e���I�"�)z���y�M6�I���)�+�RI��]|QF-�rjB锗W�n�TL5_1�����9mUf`P�;=��  �D��E!�w����v����W���Cf�e"�æRV> M
���8���7 �w!���O��gFw(ߠ����5f�je �O���^�u~:ףj}����ĤR�.���4�U�s8oa�̀�zѡZ(�4�i(�_*
ܳBaAl��3�3������wP&
YV	9������M�D$0w�A5N�r}�f������zj�08QWr/D�+y�/J�����>�(	=.��puMC�d��F�=�W��v�(
�������Ks�$jj�%����bt��х�/�.Xq"��AT m�,�T6'n<|n��m��$`�S���==�ᆮJؠ݄�3ѹ��ܫ P�ֳ��BSK������<��κ{.�o�����g��O�yb;!QWt/d*T~ܽ>�8{>c���WD��h
�����&������*�����'���?pd�$�:T�\�g�YD�Z;ՕO�ȹw�k>L��&�}A9��L�	 B>:CǱ��� �
��C\�v�n��t�v5�d��OKW_x�����A5������5���YR�e�ʘ�=Y��C�|��9�d���`���Nm��Z�ݎN�H�I���C���ߋ����A�F7\/E�yB�O��p�̽e�"�٭/6	�
1{��\-�1*�w�^�ۚ���k3��]�)|U���Kڐ�G���u^�2CQar�c��?:�����X�`�՗�
������8�x�]Jl���:˜3�ޯ��]��ٽ/.�/��EWD�>O�<@Ά41��5����ݹ�-+W������.��'��>&��}V�,y�'��bDO
\L�C�D���2N�CC�� �����C%���H�X��C��7/���ߌy�ZN�͈�c3�����[����d�h��Pt��jD���>&��ϢYY]^@�}��2��"�Ί��)���O7{n�d�K�����Ј�D�B�q{A7���'�� ����s�$T�;���PR[��ş/�y�Er0�x[(MY@�"�"`��YF%6�+3L(4:*����J������o�������n���?��כk-�u�_�G�@�:r��K��F��z#A
)?,�I���&��.�t̐&U?��%��3f���1fCI��^��|���C�e2o��t8��Q�s�~���d�"NrA�8�M��䷲�T��@�ϟ�١ �M�?�H} �z �g`��)���5�H��Q�o\�o4���B ��fr}���p�޹D���@�;�:Kb5�tُ/���ۯ!؀P����G������b��.)�K�u|k�U]A�+��iv�b��h0P�L�@�|�61�'���f���R�|\h���]�BޑI�0�EԷ4�'ߞ6=��zPti|��rkF�N�����W!x��00Z�KX�x�|��N �F�#7��Bt�ܔ�<�U���U�E�_/~��mvz�Uiw����µ��XnnD�+w��f��������]]��鱬����"��j�q"����Z�hd�5��\�#�#��ƿ�q�+*��D���.>�W7��Ð�,�k�JNdu�3�S�*=���U�i��ߠ�q����2e�K����^c��f��c[�I�w��ã��њ�j5+�p�@�c��'���ȱ�hӑ	W�X�\p
:4DQQ[��F�J�A(ʴ㡫`�`�;h�f�UZ�Cg6.m�m�ͧ3>�ٱL��l����/W�;Wapi"N	�l]p<e�!�堖bwa�ݓ9'AA$`i�ﺦ���o�v�L����Aet����|��+���Ԟ�4yyEӡ�l��6�Ax�OJ,&�6�z����	26�3G�Y���NRB~�iv�z��u��}+)n�CݓaDMu�Q�~%ᢣ��D��%}���ee���&V�}�?n� �*�/�N$�T���i+�\,�J�H�.2f�XO~�L�"	^�p�J���B�L�+�����w�O/����̎R]cF�N���}�2HT���8��x�g���:}�0���"�jͿ��˶���M���%�n{]�<$B��<�KK>�f)�Y�*��]Ӹ8��L�F��|,^�'��i0Y��a����ُ
z*i��-�a-���n���6�|���fa����C@f������Z�I�#���<����ebK�+�E��ؿ ��%�4e��[~����p)c��d>�s���l�mZ@ �)K�(:1 �%�%*���M0�4:����~�;b׍G�@��Q�us%��7�ಪ��y;?�8���>žk��>K4�~,��>���Y�ε��y ����"\�A�K�Y��r簾T"�D�d�+����?)
�T�����Y5�}��MY`^D&p�UW�_%�J8�ַ6��Xھ�#"� �:1�L>�#~QRs{�h��T�wXQֵ�@���ܰ��E�<�������r��Xdۦ�/��Q�o+3푆j��7�U�ZcΕ1y�@��i5��B���h�̂c�Qr������ձHE�X?�=S��F���;n�N�@2��Y ����o�\���8�qTzeׂ���uu?e�O�F;��Pz\-l�JQ��7� �O&1n��I���/~�z�bu��玛^�	B�W�(Hрa7&Z������k��?�c����؜x��C=c����|�	�l���ˬ�kCE��3�`ڼ,��/�}��iU��p�.���-�����z
���n�^������n�.��n�����.��CBi��w�����}����9s���;s߲y��X>��ȿط��ю���s�e����\�,T��P(e�T�ރ�Ŧ6��#���1H������Ħ���e���u����	�S��Qj��*�	�7��m�Ɠ�H�ե��^u\\IBhh�$(-�Aȵ�f�Q0$0Lu�J[Gb���e�(���Y�OX(wMy���C�FQ���<\j�ޫ�
������#��g9uM�2P\�7�$���l���&8��a%Ұ9G\i!���1��4=8<M��D�sG�R.$8�t�i��?O		���{�)5�A��!i!�+|cw
W(+:d~h���'̵���X����8)�]�H,��f9C�%�c�z���CF��"V���ĊەC~�E"�Q���j�Mi�B
����ZS1j
vn����&��YHL��y�H�R�#�5�������a��8�߉���l�~�+�YT�w�?�`��;�-�[ڨ�=��[H����M��	e<p�J���I\�V�T�IN��+�G�NPʏ3�_�6��ް��&�C��4����l�;�)$�@\=z�,x70�{�d�|��즨�<lyg�D�ж�����gBi%����&4t/��-�NH��i�~?���y����.�b&��Y]T W5���B{�zGL	���`T���{����F�Wخ�9{��Ӻ���t���|���{v�e��$M�4 }d$J3v#Bxn�C�i �pG�����p)���{��3a�_���.�|]T��5
*�I�{���@��!fo��p���>���l�C�_�Ptq�P�D�Y�`�a�Du��s�����8T� ��:�	h�����\> ��/P��l�xh��s�W.L��ў�j���ޕ_m��6���+Wb=�ڰ�l_,*u3��W��C��Ζ�q�:�M��W�c��\�>�	��q��H+N��7C&
�NR�Y�������()������
ҍ�� � X)����&#^����Azr_2��_M��!_�a>ሃ��k>������Q�Im	�imD�v.��:H/�Ɠ~�m�7�Ó�$�%��Y�o���(l����p�Ψ�1m1�����n�oG��$$�aK����&�ew�o3x���ʊ��FGX�:��2�(l�j���p�1C���4�&�P+�eZ6:{�vpw8�pD�
#���P�SQJx�����G���q���͓^�3��Eo,���s�Ϩ� K�&9J�04���yJ�h-�v@���P�����TCoͨr8��%�T��c�_W�Uz`���o����O6HW�+��Н/}!��7��5h���{ 7�'E?�v�F/���K���A�ra���(a�$fx`�ġӨ�C����Of~�䄧�DG�
�R��?i����p-u���G�C�"��/6�u�X�A��\�	����  ^����-��	T�v��
_p4�<yk3a�7ü2͜��:��섕�Ge�"�l���8"w2N��|�yb��e������g���2~�6αv?k1�~<�������ƀw#6�[�E� ��F��F �Eڂ=B�@���_p��\��^�ƫ�zDǺ!�fK"�\�^��/7e�vA��WzD�,:\�����C_#jk��F#	T�QX����汃H�̉�i��2�-��n�����%��<�����O�9+a�w'�߿G�Fي�%MH�_�:��*��UT�ڄn���Ʀ�e�x�LD0�?�E�����&��5����#zf1bqf�ۥC3�-v$/۷�ùW�~wbz�^��Y�~���|#���FX����oɺ��PYH��O��6��|���6�	�DnVW��!>"^��m�9/Xg��τ&d��*��FKD��G�Y�g��#E"� ����� �#Vٓ �=�{�h �����B~��GL�1�
����*& {��@ 4��B�����:%1�`���x!�	��k�~��:���,� �M��(B�������q
0�����c���]��L�ڈ�L3! � �7��׌��ЁvY��x���7G�$��dX�@����Ƙ���]	���2�C1�\ ى��i`僀|	��(`���`,����� ��kC`?���<��_�=��8 >��?rQ �HC�9�L�_3�L4���杋�� ���@�=���SDv1v2���Ձ��F��y���|��}�O���c�ՁG�z����{>LsMD8<D7�L7(ژ�<p%�,7���p�D����fi�@֩�7��\rB�;8�J���R��U6ǇX�6M��T��&����da\�PO�#A|A�A�m�Z};�$��	���Y�;�}J�O&gI�r%���yB$۷."�X�(�c]0�(v�"�3be�1��u\����P��T��$�Y����xu���(�ڍ,sM���X�b*>O�qGv 8x[PR]��f\�`)Pg��6���el�a�򠗭��Z�(*����g{*v�ct���$y�"Ui1j����H�"���zH�'���td��oHL�#䃴9��^&@9��~쿏�NC��RG=��Y8����$�@@��m�T���%0� ���$G�^0w+aC�#$������ט`�g$�L���Ag�t۱��06��^�����֩\�0�G���R��)ZfΘC�<(��}Z20���8��i	�9�ؖY �m�����7�~Z��x��ե
s42w��B&	��J�Y8�ޙ��:��F/nǬ�2~��ᩰ5�d50�Ӥ�2���S��W�d�zش_ْW�@�����9��Yz���G�T�ғuhm�a��+�6���wB��9����20
�A�� M]����Fa�X
@�~0I�{<�۴���)��|��-X��n,���߯�0	T�4i:���)Af�{��#�LZW���;�����z�;�K�Z��y�p��R��A�1O��GK���ɹ[ۨ��%eZX.�n%+D
O<�\��F ���?�'AKIɏ]Ϟ�w	�ƢN<Uj$�����F�C���������U2e�T"���5��+Čp��y@�k\<l!�mt����_[Y�c�Ld���B��RvN����Ǒ��m{��lbIJ��&�8�\j�2���	�|��R^0��B�'�JBNG���(�.���ç_��L <� ��b�R!qh_��yD��4)!�s�(����W�G������eպ��/<\
����,.$��W���
��ݍ�rI�u���c�Tn���4�����*7�]"�W�%ͳz�������gZE��� �P�&->B%��Q����Į����9�x��=�r�:��7��M��w*	�ˑ�g5R�uEy��tk��)���%�ؾ�˘�yғX�\+��Y��? ���N0
�)f~QH���.�	bs�_��Z��2�5ս7���V��výNr�Z��h}@S���ߋNe�q�6X?NmT����m��m����ѹ��_#�v�$�U� ��~��j_��H�\0��@��"<li��ț�l�n���AZ�QRJJy$�9F��Ht,�����H���o5��kfb���2W�'x��;�1=?�0�KN��+�����c��;sXWQ	G�"��4c�����
A�,۲خ߳W�9�Uq�W;s*�XA�,v�_M��i�2�_�/�[7��v�HKKW�yy�|Kx�+Ǿdm>�k�_��z�1�D�*Ll5�>C�Q=�"�D�emP.�X��]����qǥN�<��ieE��J^ş����vn��iU��}�g|�'�ڴ��	��\��KP= ���~�Hy���1om=��$V�㝟x�t��^b�a��&(Q;3�5X��6�d_���ǣ��S������a����@��գ�n���ބ�adm�#�|��PmP�n�f��T����TXu�y�u�U����_�&ݾ~r��\Y[/�~����Uj��ū<X&|k@6���3 v�ga�[O�xz���F��3����?�2���/��u�O%W�?������0ޫ�*A�u0>�H�1ޛ�%���OnS�qMfHH�(�$�k��w2��+��7��CDȤW'5�\���ޛ����ʩUg�įo`a�F1{�r���R�
���!O2���]�v�� ;�h���꣞��ХAX����5C��q�l(��8���j��6%@� �E�US5��M�R���	�]�]0���G9q�����)�=��G��C'��N��"�[�I�A?O%֭���2Н�����糍�_YPy����v|~7�Bf����,֯_�q�|��>�Lxh��l��Pm�,��Hx'}��W\|��r�=u������:*��<5}��Z=�;O���/�:��KU��g[���7\k$�o3e��X�_�(�\MS4�q����usg��M�nGG���%x7-_�]�O�U�Zĉ���v�X�Y4��-����@�Iŧ���w��o�Ec~�'�6V�E�wE+t[�P�##qJhj��^Sm��>�i�_�e���U���J�v���F;��%�����M겧�|���3��Mh��r65���v�g��4�4���vn��kIs���'噿�t�1�=�����2�xj�ٶѲ�M}@�L�+��	6�5�-c�f.m��f{��}F���'�򢜹r����z�F�~[��������g,U6'��S�H��l��Vos����%G$�6eH|�{{ζ(9qT�H�R]�i��b��YAަ����lXϤ�2I�NѶ���QӷQ�*:���n������0F2?��>�>�!��ԿY�Q����j��3I����֑����	_��댏���5�Ŧ�ٰ��f�@��j3�|͕���rX�0�3��������Z��*o�J��i������Pi��C9j�(8z��hT4-�J'%��O�,l�;��]�`�f�()�;�f��l]��������@j5�U8�w֢���}ޡ�<~H�	�T8]]�4|�1x[�ت�fp��
����m%(͌�R�vxr����_P�!+M�5k1��s���Ό�4���EcK�Ϙ����ٸ��R��>�m���6:б$�Z�� �Rz��7�v͍��8��p�]f�}wδ,F��@��T(^}�;�/q�j�O䝮�+���`�&��D�0*m՝�E�+4f=zH�\�,1e΢qG���st~^	C1�;�q���'������e#[��ơ�w�J֩�����m�p�Y�~Z�¢��O�5*�Ҷi���b�39n��\��]2!�I"��g��q�����?Ȉ Y���&�/q[1���ϣfM7��>=%�w����]����x�5d�`�3�AtC���﫷kMM�hGɑ,z�2W�辣>��!�^��*�[���&
A2�z}[HM�]�I��������h��ao��|��՛��aC�F8�����dɈ�
u=ej]&!/��I�~j~ɬ�m,�f�B�̇�8ң��Y�6<��7/�ۭZ��v`Nc�����yQ��Q`@�ڵ~G
���e,a����O���2����D�*��4���,Xw�z#_�s���ڝ��v��;=�ӶF6��-��ua+C_�� j�'6[�z���S����~�M�'���cg�Cxwoh��P���x�&S��U�\��7��Ļ�����6{��q,%�Z)���j�C1�y��&��T��&	�M��F^�r;m%��jg�O�@��D�8^7]�~�¯�������_}f]�����)XF�p�U-V+.�d�U���6�{L�WC����8��N���w;t�v�m>��s��WV�|�>�y�m�N��Hr�1��߫9`�S���U�d#��C6d25�a���`禡Jq�[��T�f�;��]WǨi���+�a��ɡ�'YY8)c����r�R�ۉyh����=���_o3bͻ�KI�#��ݿ�g����?�Y��t.n����N���0n��[\G����UC�ۄ� ���z�".&,N�"�2&%K�ޖ���G��p\O�g��흴׾�E�@�<R�վ���Iemd[�������mY1,y&<Q�{%l|�t��V����G��F����5�l7����H�7�J�GsӶC���lDkd�q��y_@���T���?b������g1D�~��6Xq�vV5�aI΃���c�������C�d��n�n➦��n�Wn�K��;���^���ܤ�9�㜏}qK.��y������x��b��j
���J�Y	����[�ͭ�2�>�BR�)��Kҋv���B$����I�k��� %����?�qЕ���^'YӘӾ�@e�KN?�#]���ڨ��R��'����ϵL��f���J�7����ܙ�Ÿ� wL�P�7� �{��C$
yLGP��1 }��

ڈF� �/
5�Y����R�j��
���EI��;��x�'̵�xO�W_5��@�K��ymn������z&ju���-�/�Y�<|TK�3.7J���Ê�Y�$���UJ������]���ى�Q�I�+�1��o�I�p�rz�Dj�n߁�����RPk��ت'x�+�\���fo�gG������[vxʴ�O�Jc��!΃��Eu����K�ndUrR�
��Y����C�h�#����樓c��ܻ�@R��%pzn/Fܶ����=�=7��� ���!�����dU��s#�=�aA�~�הå���
��_�9'�TM��vfڲH�#���\ҶŲ��gB ������
�XP�[I>����]�E~�v����;�315)�YY�R�C���x��?���a�Μ�Z����go`��TЦ"E;c}k����p��A��5�1�Q!�Di�B�u�op�8}��=^����uO*�����{.���8��$+��{?[�]��s톇o%L�ޔW��P��"a�����)-�B���]l��V|Lq�{⟤�g��V~+>=���o6:4��t
��T(������[��R{R�8��ɻ�5OZ�8f�r��7��d�W��xb�H,4���84]��ܷ�䐃!�=;�����	^o�FL�#�5xE��x!����m������]�����IGo���s���%���n�*z�F������qo��NDG� 1BG<z�skA)N���i/%�oy����:ُf�Q�׿���2Jw��m[���J>��uD9l�F��X�ٸD���I�)j�D����C��#!�_������zؖ��HB�*Z>{��9È=��A��8/j�jc�؝���H����c��,��P���A��g��j�v��
)�l,�����+&(h~��~w�����:X\�J|�$���N�l���d*�����9iV�$q�i�⓪9)�&ڵ��9�	�ߖ+�,�4�J�4,�^��u��sf~!��o{54�ƣ�dMv>�R�$�����a�@~3�A#g�Ol-�l�~�R�Xe�3I�x���s����@�M�\8�(�:���&hH������X��<��PR*`���ӧ({ *|;S�H�H#�X�7�	_ ���mS)�-�m��āg���b�"k���g��3㧣S0�m��j8���F��~Z�h�Ż���fC��3�ë�E�$���������fo.+�'s#�ȉΥ�Ѳ#�%n9���X����2#�S�O����s=�|�j���7q&$�F��6�����w�8(�;�e���e�Z���@�r)�oo�Mrko7�g�Na����_��!�G~7��{��F(�\��or�|��z�p�Ug�T��Pdq�ט˲��e�����u~��Q��ޫ{w�G|��@w�
8L��x�����B���Ƿ�͹Zt��mu�+�_6����eĄT�4��Y(�YNpHX0�\��d��N��\��"��qk�b�n������ڈ�x����/Ls�z4"x��_�Y��D�n����aj��.����Gb��(����L�["�v��c���G��K6��!H�*FIs�������������W��Dl��1 DT�����L��z�T��=_K<,Fg�e ��
�d�td3���y���W&��|��0����o���9�YǙ�fC�ȇ��-�Û"P��NG+�O�\�u�O-@*�r�v�"�⃃;de>r�k��q�i1��jI[W���(b��xE�Zf��l�g�??;zFR��'n��pt�y�z�O��=k�AGl�U)���]'X���8Q_0}g��%����n?��:c��$Fw{X���{��یVDn���)fw�>�]��;��3��Z؝W�.��I�OɋB��M	�u��:ݖ����:.��!�MBP�]P;DI��y�ʫA؛�!I�G(*��4�ȷ�2nn6�P��P����堁Gp"&f�E� �������oE��g��9U����0�����������%� �i�ȕ� dR�p0<U�/Oi���P41�����5�7[���SL©7k؀ur��Vq��h�����e���,'C$�
�qC�?>m�T�)�`
��P���fٽMsa�Y��Fq/p��Q�չ�\P�I7�@�!�#�,�Z������|�BZ�r�M}�FΞ��{Td'��!�ԙҝk!�j3��>8Q�	Bw�nq����#��v��yjpؑq �h$]/ �L	�RЛ�M���]a�c�766��-Q��#$�]Ӳ�כ���:��O�D�*=���(lU-Z��f��P�:#����6���
����w�Y�W�f������Ê��8 ��5�ݜ[���~y�&q��  ��m�P��q�R~&��/�p ��/Z�����]�4�Q�TD. ?��~jU_ۚe�gi��ݮ�Z$j�hh`~��rkG�4d�	�)n
���-��모 �w�t�r&�gqo��<�p0d��q�S��i!��g@��	/~ՓRٺ�����f���fz��$л�m�
���|�9Aշ���OO�7�O;/&�NO'��[�c��j�����ȧJ͆�Y݌iU���:WR%^����`t?����vW���@�9{׀ϥ7����~�r؛w9L$h�C���.G�Զ��翃8�t��WT��;���ά昖�Q�a�4Й?K��lji���&�vS8`��$]�^�������/�k��}Mޯ�+�}}x`6�y��]��śY�L���
y�b�4H"=wL#yq��-�����zI�����w��)j(`^%^YM�;��k?H�#`�h^ȴ��z�Q�mL6�!�ޮ�x�6���~5���n�o�>���d-WQ��@?��[��2ş�o.��c�vB�J�k���Q����g�����3Y ��&��!���+�¦⽑1!C�2�؈ٿH!�ԄQ�Q�)���&t$�q;\�Hrl�B��\��J}X�B%2�>�H.^�������M�ڃ��Pb�2��V�ـ��fYԆ�u�]�냮C"B���N�8Q�!iTu)
r�1�Ȃ���%���`�"��V��}YP�H.�ʗ��7R?�=Φ�����^~)@���)�i��	H��moy�;aW�Ν�l@�t��`H�����5�����"2$�']JE�!�c]�.���zs,ܷ-��(X�nr��+ Y��A�M MQ0�6xYM���r�5���7�3�Pfn�=��T��y1��.�7��d�:@�{h|������8O���g#ٟ]�╡&;�x�v�-���[��)��B��gRj_ޜ�i�^!/-`	���h�вe�j��J&A���3XE��%Ƈal@��H8�6��t�YJ����Y��b�f(���,{�ό�t�)���x���:�����y-�%cz��n/2J
��2���l���4�g���$�,���a�J�G���Mޔui\f�����������?�a�����97&gi:Z=՜#��
_��]�;m��ځ�[����_�V�$.k� r?����srw8���ڲb^㊚tɋ�� ��qj�^l�yڒ���>��P:J���Yo�l�?��}1^�f�s�����;��w�� �W��*��W����ï`���m�C�����j�-_�?԰a9��@������N��i#ˁӄ�.��l[�g�^��:�n/���$έ�(hJ6n��؈��v�5a}��&"�g��9Q������)N��y#��:�y���Ȫ�����z��{����fUT���l�����:���獉x�{L�ʴ�d̔��On�c���Z7���s��N��r�	��Yǆ7�pȟP�o��-S�Y��>
���Y����& w�5�Z�~qI6|�6ے��ъR'f�1�ϊB�~R}�v!3�����N�?_o|xIm
p�0!��$���	�g�\0@S(L���1	�s�{�`B��-��^�s5��GK��f�Am���+>�?{\�d:����ل}�78�E�X<B�H�U����0yE@JJZ�٬�#�̌�M���(����P������yO��y��oK�l��2�˦5�"��b�L� ���ojh�uk߭fu�Ƣ�4������J�U�k�珙�Z��M�\Q�z-6D���za�:��W�>���N�8�_a�[�����uhE�d����m �q6-��P����'�F>1m/���?���;�b�i�fy�ۀ������^�(f�� ��{��n2������0%ox]�̙�]�ޏg��`�yv�O��~�̟k��@�|�z�.9����2���U�w버�vۚF����q������+j7+Q�-`=<�:q����7�SXpd>>�H>n�Ds�
��*�}inv=�GVB~x�I�K5L��,(e�%Ԓ`X7W�*�x���ԗ�`G^���u�J�Ro�Y�H*�.�")��k�۽Wm��Z���/�vI���-o��4���ޛ��_W2Rn�E��� ��sv�����/^E-��rȅ\��4V�s���u$�q���>~���8z�[hr2V�E�]�U��N�l��癭$��c-v�R�/���Uhl��y)bxnW�n��e.���`��L@���{'���+�T��zye���:�LT�J\��]^6�&D5��
q��?*�w�R4�WmY�o��oߟ���A� �n����M^�-���7nhw!u��
�4��7"���V{x�u�����#B����1c��G�e���+�\���!�8�.�˨�����d��֦,�j��j��>d|��1�$�T������b6����k�(u0,(�/	�MB��N����T3���h�u�CB�g�˞9�B�'K��l9N�$�M����b������Z�ga���*��b�HH��4��@gͧ�ݏ��n^Ϋ$�%~��U�Ȁ�����X�4�i6?B(��Zu�8��Rw��'#��߆�L��Y�i�閍;QR�6s|�)́9$� ��B��q<_��#��|a\�#����Q	\$N��=j^����H��z�Mrˀ�y�Z�V�C��QeU�2�Sz���#"���s��i�2;�e�w��e�^��">�8h�62�̅�%X�?޼�V��Q�=]i��]o�=�S�gI�/c�oX�q"Ǻ�mr.�/�rq���>�s�ػ[9�_���)[m�rg^bURiE�Km)r�S�Jn�9f:*!2HÆyf�N�S8�X;��j�)]e�S��Hz���g�[^t�#X�tq�9�Y�q�p�s�����U��y��J2�n`j����c5e"�"�n`����>�R�����\��tg-&QՋ�6��V|����������t�b4Z�f���$�����"<8���8E�$���0�l�mڧ�#|b�*>qV/�����f����J�u���.�����D�<�7$�D��<��t6�+���T�9�8�6�'�������"�f�ń|ؿ�,ȷz'�Ũ��3#�����k"��b�%���xN����n��-�lL��&�[fg)Q��K�4tBc�ִ���{B,��5O���͟��X�6��U�-�����<������ރ,m��I4(�GX����󡤊d�-t�8&
W�o�M�y΂B_Ү��.dYZSd���d�׵����rF(3o7�����WS��x���O/˚X��ұ3�����TA��B�u�?��>�]��(0$�y:l>�	*(���v�a�t$�v}B� ��x�!�v�΀��Nm�w�7�={�}���v�n�m�	�#r#�y��`P���}&���Ԭ/����u!,HRlX?�y�h|��\�h�1�w�֍!EAN"uv���]��C�y��$r�~0z:G���<nD���|n$�CՋ�&�r�Nԝ���8��yP4��<A�❎_W苾��7��Ⱦ�����?c���gz|j���ɲ����!D�d-���.�hF��x7�󡯹GJ84uF�ɥM)Lbj�-!�B�ǈ��8V�ܿ��%3���=6�O��x3�⵿D��ў/�1�Agd�EDm�8�f�/�޾����OE5��o�}�adv�ԗ�斾��'�D�v�VɴH�"��"-��s�kܘ~x����X�#�"}d.Y�;Dx󼤕m�-�_�n�GK��x��������߶��&H�{{�4�k�j4�pr�Է�-A��>����{������oÜ���x�G��2c1����p��4�]Ь����`��]T���z��~�fQg�(e�x6�M��I�=hgH(�]�'�?f���=.�[�H�g��/�h�)�,�|1I�6�d	L��!�zt�������@��Mh��ʟc��ҵ�m[�s�SH����|��f� q�d�pU�~�w�r����w3�e��YI��R�r�=ٱDH���kC��Fl��y�w���3]���B`M�����h���#�E��H������n8��`퐲
�K�n�EU��5ii\0�$��%�Md��Ekl���!<�E��1��[޻�iB�)�e�t�}�������{S�@��0��0�d�yQj�S���䟃01��m�K��U)\sB��ŦMxBG0�1
H���&J	>�q�f[P�f1���@1QrX��2����գ��Q��O�D���s\���L!j5'�Y�D`����g� �0�8l;��
"��96�)�A�x2d:)Da��R�,c�{Q���JJJ�@�',E�$��̚$P�c��t�^��T�2�%%���c �B�sCxE7�?1������YD#PL���|���>���͠% ��'�GH!z$A��_�L \F��@q	�Å��B��,���i$�OC�� ��A l��DY��� ��1dL=v�)UȘ�a�7�Gm�cF�멂B�2&��y���<d��;��� hMA�cԐ��@O~@$���(�_ � # �2?��	� \ ��Lq�z�\l���	��-�ƀ���`˷@hH���ɮ�TK A����_�V����d���qBHH�����^�
Ї�	�U�7��� �4B�O|e���} nVA�G]".7B�&� n8E�`��-NY��9�"ȍR�jV�Y�X04�/
w�B0��C���� W��}k}���G.LKu������J��ݚJZ����\�Aue�\D;j���ҍ�n,}�He��
�su]P�����R�֒�y�z����K4D; f�hp2f�U���n�J(��t���!�ȡ�ЬGXE���a<��|>kŏW���%�Wt 8Z�� =J"�%�ݖe
�֢ʐ������@�]��z�p�}�9W�<�II{���eL�:p�)�Yc�z�)o8�PL+顇���>�ô���j���������3<�0�1X�#=��q� <���ML+�����a����ĢD�oH��F���u=���@�A���ւ�B%����p��С�N_��Q��ç~���MAe)z\H�T�Ѫ�|W��LA�2h�ܲAl0���;1�nO��%������z�0����RZ���C�d�Jf�O�[5�����.y� 0�̓������. u�OH���ej����#��J�<w��&%>X"њ�{��f�.�%A��H�׃5&$�2M�K���	M�
�#��Ats�Ε������=Е:�+�E�"D@�����YDm�����u�"}�~nyv�VZ1� �$�VLF&�2�R�6</�Ĺ��?�CaN'��}G�̈́����CH+�m�+�X�9����`��\I-���n�C?���B��p��s��Fɰ��'��������ԗ{��=��j�Ik��%3J�mw�]I�bO6���C�V��&B�� Z0��6{���|c$�4%l���=#�2	�9�F@]#,KQ4a��A�[�����x�;��Sk���䖂�Z�T5�u����[)"��2v��wA����[����?P`3J(㨈H%99Bz_��\����b�,�v"L?��D(L]$T��^H��0�a(�55�0����J�JN�8Jəz�!���Mͺ�Q�!۫u�4?�k�� F�%,���,	���/8})N�o2Wc�eպ��̷o�۪)�NK�wte������d����3��R@�i�:ޝ���z�TdrX��Z(�Bd��g��	���P޸=�:`�Y_0�!BOa��X��Hsr�z�)�u
,��(0/-)�v�z|�v��]d1�ߥg�i������ć�דɝ�
tb뜾�%�v���<����zT���PW}	�3�,�{hx/�=��$D�׼�<�z$"�Ӫ��.��`.����2�&���K���C���Nw�2�m�J+_n�%
dͽ��J�φ�)y1g�������:�m"�b'�L�pU҄���@���7��w8�� �0`P��(�����m,����>sl��;�ii�Hʭk�FKNr80ڜ3`�;{�E��s���i9��~^آ�GC9p�?�r7���#�
���I��K�i~[��4,�����0��`9}`���c���eE?�a9O#W�Y� =�f��с�-U������M��@��z�G������8���.F�?$ӿs�C�/��ԉ�6�j@�V[;�����	�A/(�O)/�B޻��+0'��u%8lG�`70vk}G
͂gi�%=��B^q<Yn�����'\Ee���םߴ�:�ۜ ������.C�^ڣ��k�tf�B���<s�n�W������ܻ[��n�͏c(�\푩{��]��zm�ٷ�6W��w{�y:���УPJJ. �����RV�g���У����̛�O�]CԳ"�vO��?���`�� �3=%I����@ޭ�D�uE&�����o\?W��=�ʳ���My�z��3����4K���g_ֿ=t��i��7��j��
v���������w��0����F�Ni9V�N�ibF7	��h�=[��~��M��z�tzZwv�����Q���dK�z(�l"`<p3�+�y2��_Z�����e�&j� �"�t�9W�\c�c���"��-�Xi�F��Vp_ֳ�\��rdL�r����;.��7�0S'�DO��E.
���EW���zsa\�����OnE��J�*#
�*8���B���DU�Ye�[Rum�FS�v;�Ы��
s۽�|�^��/�YIH+1]���5���Un'�+_/��U�	������|�K��rr��Vh1��VQ�f�D�Ƶo�6�x[︓�x��#"��5o����ѓ4��I�(�	lc�|&�����x���m�׹���c���S��8ΟK���{C�^iԹ��\a�����WN`��<|���&}��ix��(_}��*%}w�\ܳ��'X�J�h��R^�:�k�뼞�E����wk�ظU���x7��sy#�	]4.�V��t�G&�?0���㥿�7�;�8��R}<�(�&��;BMh(��A�K\Ҍ�x��B�:�5����d3Ld��U����w	^��H���>^v�v'i�}q"�sSl���Q�����t戻`��
+�����㺂��j��Dna�ͪ��D$Y�l�E�o(\&���a�\�?CJ���	+*��頱7�"~<|��:���o�'x�ƭ��ة���>?P�i�V��9��uP��ww5l ���6��"��1�r���Ź�����3�R��V��u}
��<&²(\@K�_L�>��2�I\wҶj�Ĺ�J
��#탡gSBjF�ƒ��
k���#���7�x�����FOQ���g
�?���:ck4��������Fz��o)�1;-;���*�[��?5 ���Mit\d���Ģ⇗�д��_<��+Q�ZQ64��Mւ��e�R��W�*���?^�^��DP�E",�̭.��u;���R�U��
?F�AVn4u?f�����^������>�P�_F���/��q�d�m�4�,��h��{qy�˾y�h�IP�?m~J|"y;p��$�R���F2�h���%��ػ�}����-EG� �E?��l�	���M�C��΄,yL��4�g���}��5�8�?C��.��p��٫4�mQW��,��
=	�һ6�e��H���x,g�:���.fs��@J�(���8\ǷĆT`h��n����t�w��f]��6��@�������$��,����}I,����j���66�P���k]{i�y�oI\��*&��Hd�O�Q�:&�D������7���YC(R���
Fwy���1=v4V�|˪����������i֋�Cpw'wנ	��N� ��[p]48�eC�8���w�9��StwuM�SO�T�HHĊ�IdE@H�Y,��[\�� ��o1�x�U�AxÜ$��i�݂V�%��SC�	"`t��e���9�D�x����!��F�d�������8smK�XWE����5Ua��i��Q��K�4���x��qS�Y�q󩡀�XP��Z�V>`]@}��Dx��D��v� ��l4P(po�o� �x�6ɁE�����{y�<jZ����mxR�-n����������*�rg��(��V�y^(<q���J��h��u[�,��V��ŗ_(=�hv�d���r����7�%0rW\�~��72jʱX�f� ����].*�m�2Э߉���s����:�����3��<W�#dsDX��⌬(Y}�[�6,xb�NM�%�̻첎���jyJ�]�2�iw��|l�hx�\�s�ò��b��45��9�*�p7ћ�yR��U衭��C��<&5_��)�	��x���rb���{s^�u��Y�ga�F�u[*Cr!�r��� h'tK��R*H��go�t��V�E�z�ѓF��=�7�w�R���o�UٌzL^�?��K��(n���;:�\i�4"t-�4x5֑_|��MX<�׿`Մ�}�G{"�r˶��������z��2q�^���?��f���|��G���Sr�s��&_����d�Z��2�_��]� &��w*Z�r%[s���a��(}�Z��gVF˦I��ܲ:���#�Z'>����dv�w�)��]��	�)tb�<+Րe�=�vվI���妎b���H�<v�7����/�z<:Q�?�q��M:]����u���ʴ�T��΅MR �<2v�/�J�@8��]D:�Q��%2gh�:}�,�i��9���o�/!�dwYV���^q�
�Ԋ-�m�&dl��r����뉤�*�U��6�b�M��]�y�1=�$�b����t�w��I��c�ȤR�C_�`_�ٖ�O�=yqa?޵��)�q��9����6X�|,ϸ�'0X2ϴ��H��2{�V���(��3$��s�*��/�q��#U?��@�ɋՃs�'C��/}�6���{��F�G�ۏ�\���i֡�Xb��{H����|���k%}�֝,7��`��-dI�-z'�8�:am���zE�Ǥ1�hڹ4'\7���+U^}�j�r��@*$����n$P�N�-�!p�ϩ®��l����r�Ѡ��r���@?�C�x�C{��v��K"��^G��N�WN݀�������51H�K��K�����e\i�NǺC o;�/�d�u����%/������(�r;��`���//���c�A1J��/n��P#."��h��~�H��"N4\veÆZl̘���!�� m�4,��K�j�G�iR!����۫=�'u�`'��&kt])mM�Fz��9��'W:�OB5?�����ƿ���ǘ��3.����������n*q|ij�fp�w#��*NC$�v��g�>�i�����_��<xT�t ��<K%�6��&�ƥ>FW�9 ѢЋ"�f�|Vwx�ơa�h��j����l`����[u5�<�R{3�-+������!�����)J/}���02.� �4���m��h��ލ���J�|Q�aw3�u�K���ɠ��\��կ� ّxPIG�PF�U�jd�,��rļ|��C?��í�צ�i��H����+p�џ̂�����#+T�
��N�z_���U/���#,��dQ��@��Kd��Ih��8�	��
��#w���2���H���x􍖟u�9BPCC4u����ۡ���B����1����n�{�Ȋ} �J ��L��eE�'RȖh"�/˙@owp�=��[��c]V����휾�V�R*���~��Y��S�]v��k;���e��*z��h�̞7�!&���X�Y^�	u��KP_�Y��0P�7@z��$�oC8���ғz&7RW=� �F|ƾ@�\>zq7q�J�b�dtՌ��](K�m/�����G!Z��U|�.�>��(}��~����
�)wp3H�2l��F����x>T�����5�<DJliYm�So�̭H�" ۦ:�j��t$�a���$V�Q'������|8���5���$����g����m���W3�XBlы;���O�庋�(C��H ���"�;�8������{ON�Y{��v�{�ͨ�
��P9)a �B"aO;%6ؾF�I���ʷ,�.s[��ǚBb2Q_�J �����[&���-�?=JP�/Z����o4��~_�(/����;b�L�U����I�ʝ"R�{"��d� �'ר��� �V���[e*W|P�eQ�ѩDve ��>=�!���m1��bd%R���a�����(�_ZI���?qб1E�d�.���Q��Z캨o�`NQ�NX���)A�l�w"H�Z���b��A�[��k���n�Z-��|4��
���,h��h3���&�j��|�������o��@Y�RqH�2葺�����}��`�c��-տ�Ge�n:�H����e��"�V�%J:J��B�=��i6�*"�7B�ą������6bg�6D��.��*rn��!��Х;bI!Գ�����B�X��jK3ʊ@���O,�)��/}(�7

��,�6�Za��Ҷ��7�E٭����k��Gm@\tZT�_���%F���┯��^%w�'��B���2�g�!�3���[Y5���a(1`��Ƕ��~`�uG�@���Q7!Ͻ���g"+z������F����I�?����T�P^B�G�A�W�����9����~��DcΩqB�O��z�w&:ss�d� ®z�t��3����Rm�ҽ��w�����nr��hy�"2B��Ӷ���ِtRR�mv�+�tY'�_=7L;�	vh��N��!��+�:X��'A���;���..�W(�j�5�Z1c��t��v�%�p�Ә�M��#��\@�|���/rW'��f�F,�[{�Ȳ�~���r����6Q�x윗�(�KPV�;TbJ�<$��jW�]X ֈ7�X��������,�R?N%C����E�`R
�܌���ju��	� �i�;Mo
V[�j�C��DS�@�+D �9�꿛�eN��n���q��_sI1�4+8����\��t
�x~��hyd���3�L�wE�l� S�1#q��"��������P�bd=���Q��;N1(�-�2_����b:
47��v[�;\��b�^��&�*;6]��{k^z�qл���]������{P��ǥ4)J�w܇�TS8&�ʴ����e*_O����4�N���΀%+�7z�)J��Y�ĨP �Q�X�����Y�7�c�\5d/�&9z_��b���	�of��p�O���O�9)�Id���1����(��{�ח#E��Of)F_.?���t�҅�c�"�t��{B�H�q�[�4+"#E��;���h�l-Ռ뚮��o�sM%ay�Q	�O_�~�oƄZ�
]!����!��[��z�*o�m�z����0��hL��V���_�yU9 D���ߧ�_�Ї׍���ޜL��Gα�[�>�˲o��HyC}�k}5��zuB!����rQ_�AR�wOY�26}�;�B�c)��������K,��0�3�̇���>�=��h��t�s�A����,	�u�<e"�l8��*����rP@�ظL*�y�X�,P}��mCF��^R�Y���x�j]��x>ˇ��wn%��l�ޛ�bq�4�[�����Z����~~*ri����{�7|�!�~�)�m~(���6��]�eHS�S� 4�-6�����V�E����.����5�+r��R~���1�9��lF�(Q�1��?��J� �IF�tJ�O�Jz�oO�ǡ�c7���r��P��B*��60�v��86��*`�J(�����T��y�S��@��y�m%As�i#��>��\�84z���:��ڷ̯�[����R����U�Uk+���ͫ��,`�g�"!/rF��.�u#���DYY^�?��ӱ�K�?k�� 4�D�=J�_���+�|Cy��{D9D�?��-���tQΗ���É�1������LQ�%z�K���OTWW_��tM�8�"��T��^{ۘ���ϥ�p�j���[D��y��@�_!HD=�B�ᯁ�)t��_C�V<��V{��dr�H�q���vλ<	~����epK�t0��INN/�Ȓ�{�7{d(b�}�]e��;��(�33��j�(�~2�����V�f�+rk�ާ7�'+2�����b�Ic��R..G��y�ngG"XKR75�p�ku�����&(��qSJW����ɚ�1M���Z�	���'X����{o��ߔm2�$��B��F������o_�A����x/���˟3�䥧Ӊ�>��r���@gBkΐ&���,�d~,&+xP<�5�ʹx�n������p�i܀�X�n���Yz�K')�(U0�����\�J����_�J=�Ʉ,їǕ�#�J"�N]j���L�����|����?Zdu�H*�U��{[8y`V�~
����a�y�Ƕ��(H;9�7�堣����YH�� .� ������S����ղi�W|O�8F���_l!���U�L ���b��i���b[_���Ͷtʻ�R������B%(�mn��I����c��ؚ�[,EZ����cf�>��SRRr�U�.�3q�'E>ί��=���U0��J}"��x�U\�?T�A�M��j׌����o7ye��q|�n�ئR�6��[[�|k�>���}��_�5�K�N�u�v���\V�'W)��5�x+�����^�L����:v~~�$�c�+����B�]�l�mN��}+u�wm"�n��b���qy�Gy!��o���Џ���Շ3p��8�@ɯ*P��q�@2,����f�-�݌u�� ���O���X�`]V��n��O�\��A��c�ҴV�1p��_�/G������xq��`҉��"'1J��r�~��D��C����B���)Uq!�


��?�X2����$z���^�o��"@���Z�/�>lhH"�Y��Y���x6"�y����v�W������'fi���g��m�<��S�8��7�̕�dv;/��c�����}�E6�'�@)�Uw=�;c�*�&��2����� 
��A;�nLʆ��`
�ϛh�������$TT�g�+'�*7�P�H�3����E�<0�#�'B"����=��sN4��fah�Og� ��/����c����:�;��綵�m(��梸wz����Mπ�Q��������������+rr"@��5����ɏ�b���e>����Nc����!	g�2m�:������"�J?�g�%�`�x!�A�÷821s-W��y���>Ƴ'��&�=]�:��f������'hb�l2x�FSs~x��$��V����&W:�֙$��~�E����#q��bv����x����Q>c��m69k�;?z�ld��,ž{~�L���C��)J/�v��a9]�Y��§*m�!u�z0TI$/����!����廁���"8�ը���;�$r�/�!�L��i�8҄�v�Z�!�XKk	�(���"y
l�4�����t��)J����X��P�"xo�iD��͸���h����djf����C9�.����3�}��c��j67�OJ �Z9�!	�H��,X��R������]0A�͙sjt}
K�b���L::\I�4$�*�ڒrwԛA�X�OX��z��Uâ���L9��Li^��Gg	��f�M������XŹ����CJ��ě	6Ĵ�	|:��;���� �c�oht1r����Gw�;��z�+�\�l��H$ܦ�ʬ$H6����<��Y�F�i�+{x������q�5��-�:��>M�J��	�'���Qw�"d�J_��&�����p*�6����u����W�{���)ծ�x9�-Q��U��m��o�k��#�\7]J2��hD�eD�����?��ֽ���C��X�������.���:�;l��}�dU2Ǉ[��oRA��;����\")��`��%4�B�;-�mΙw+Y��B��ze��\�p������H�c+�M���l�u"��Ȼ����w-���N�K��d�_�}k�Ά,!c��`�Q�V�KM�	g�]�.���~�^h��7V����n��z�馁f:�8���v���Z�Owr��{d{�J����Mƕ�G5�����6�s#�U����D�������8�k��8&�p�KWzcޔ�f/��\*[*.ʺԅF6U���ɛ�]�7���u�VD4
O��3���0v�]dh�g�|B׍D�c&�pv�M��đ�u��8@\A��Mb��S$Q��th��AJk���b�E�{�5�2�]����0DZ7�|������z���ߏ(�¶r�D�7��!0���F.���bs�8A��#ѯ��_��
�x��p&V��0�ND"QD���N#�ۏZ"�ʋL(ڷՏ9!V������$�@�q�<bһ�.�_�;R�l�$n���Է��qbuqq�`|z>��a/"��$�p{��#�1H���?��mp}��������v84 ��u5˚�OSiG]����_��eR��;��Y�X0oM��*�6>�U;�뷁��e��b��J���-�k�Zڶ Y,^y���ɫ�A��yL� ���_�߮��vbu;t��,�ݬN}Y������K���ak]�F����fj�A��Q��Nv?�ޓ���_(캗_��+��dmt��b����)>�~�$.r輫*��z]݉������)aˉ�X�)Z�ɣ�s�dc��E��5è�\��?QVģ<��-%�RsM��*^ybȸ9e��U�ü6W�c�D�w������<c���ڄ�$T��������s��C��!�� O�7�y�(m������ZX9k�>���v~�P<:�Vz�B��Z6�r�ȍ��~1". U�M�d19�l���\l7�KRn;�:�f����O'��9%:�&=�;[Y��vd��{n��~$®���x;	s���7q`��؉V��0Q�m�gu�^���?1�5h�ʢa�_��։�Ly�9;ǰ���!����i���^}h�pq2,m"�ɮ7���+������Epں�e�"܀��j{�PC���J>�oz�0X��]8������R�|J��n+r4��F��b>�qgk���k����Ã���@�|�Lx�PB
�wv�iQ�F&D�!p����L��t��U��i�U~h,'@���4��)�x�A�G��E������UV�{9җ��H�~����u�$@ko14�!jY_a�p��ZI*l!־�D��ؠ/f��� �Wg�V"���`�/��j�kz��`�a���
�G�s0p���'â�řR��o"�{��I��)�؇ u�_�Vt=c���?��2߂1��F�D�;&$C���䴻B���(�9�n&)�xs�#9�����?{Oh="_`9f��{"�=E򕇝)g	&������q�|[���{B�wo�/��2�Tžz���< �VF�$�5�.��a|�%e�q�,��Б�i�iB��Z6���5(YKV�����U�׹(À��,�xP+���Z	�q��g���d���T��T2��� �P��X�Tl�Qh�S��%l#�vZ
�u��h*�Jb��X��i~�T��)��G�����{��ϗ�Ϻ#�3�y��*V�ޮo>��T?�p�;��B�q�U�)Y*����9A�����	Ů(dL|��Sr�[���A�G�⛀��&�/���7:��	�*�34��G��*��L�d2���dɘ��p|���ld����Z��{��i�e,���C�2��@<"2T���/XA-_IB"]��k:	��,��)L�&��
�`�$FF2r60\ƄΓ��Kg�O"c_5D�� T��,�ʩu��*Б���E���h,蚜��yp�Xa
1�І�(^:l�f�J�0�L� b��"0�%L9o9 ]1��	��}�9���
tM]蚭�yBp�Ԡ���������[�	���*�Ua�:ѯ���F��D���7�-t�tm��C}`Cx�5�`��-j�E%��HǀjD�Hf�\آY�2��U�#��g�NK�CǦ�G��( f"Oؚ��#qÄv0!t���1��U
�֚*4D��/�*ĀY^U��Y�(��ǍT��b�B k5.\�'845��kvLv��W>����}���Մ�°Vl\NN���x�̆�!Z{�86�Pl,)�e9><��"�"h���p��#D�>��/���uR���Lv��?�Ċm�ɚ�,��JDφ�;���~+��=:>��_���N�*���?T*Ygr}?i��{�E��vme�:T�L��Ǝ/��a��U	��?������P��k��h�P�8T����Ăr>��b��p�T4N�"Ƥ�q~��7Xj%��Hx��%�퐙@�՚k������'vBK�R��6{\��I��q�H�lh�=xı��E4M�+䉛4�,yÝ�
n�#{��"�1��ό�9R)�\��X �j>��i�F0.��9�$J�S:�m��.��n�)�@�}�N�\�ԗV��J1��	)�N ����:K ���s�	]~��/�Jk7�t*�<�
!RBQܲ ��uvb �����;����OLF")�S�M��$��U�,=(�i�_�`�%W�+� �سy���Xٚ~{~�,�vI�<�=@�.⊆	��)���ЯLC�~qi��ǡ�C ����p�K��i���W�)��;���<��8['����C��%t��N-��zMm#��϶Q��MH��2��T<�α�И��Hs�}�	;8q9w�~����ާ<v�����QW�@(�N�w�<M�	Z@����!��l�_�@ri2x(��H�L��ڨ�$$[/��cg��	=��'| �͗����]���8�}�d���y���&>�!F�)�NN'Ԟ ��î��G�R�~�z֘"N:6���6>X�����v�:}
K��������*�D��Bʙƞ�^_��Cz�>�q~���䙄�^��>�ʵ�_Ez� ���z� �P?,2�{O�_혭������70���	7���ށͲ	ox(��;~�� �ꨥ�FQ$Ik��9�~�Җ����% ���;(�a=�Ҽ��0�ɍ�M�����u�[x��<f��])(~�rM*Ǹ�W�2M@��S�G���}P�L�o�+,w%�mu�^
�:c�4��ဏ�?tx�P�J0�v�_v�GD��;���7�x̎]�=�=�>H���[ͺJ�m��
Q��e`!�|�쌍W��H���F��B8�n�Ф�74+m�Y,�'}Z�70
$�6��O�C[�ͤ��r<���A����]�o�9��m��՘'����4�5$j�<�JE��c[J5�M9�oId~b Q���QE�֜]̈́�~-��o��\T]�6�1͕Z[q�b�$�"�=�rw�%"o��P�d]=�עr�~jv]7�i��3Ncr�ӡ&`?2��;�d����h��*W M��a�,Ǩ��om-� �m]��N�!� ;��=��£ܮP�h���� x�p��b�߁��j+��C��+�	�{nP�}(?�Wc��(�e�ɈEL��~��C����1����v��Sf��;u,x��Q?�/�]Q��r�GFPEQ��4R�	5"��	��-�?5TlP������#�G`A�|� 1��P?�w��&o�����@��4�&�5��w����d���K���7�]r��C��?n��w@y=mN'�`o�F��I2ॺv��d�ȁ�O-��\�!,`�GΆ
��v2�㈡�@KE��F���J(B[�\>cTi�R7PR�M��b�U1��bj
]..+�o���Ϸe�W�����z�?YA�Q��i۱��E.�\���1�����G5�+��f$��p�������m�b�����:'���~%%0�Gc��m'|���?W�BL��ʥ����9�v��;�l]���q޷������~�ތ?NO���V�Cى�|�{Z#�e�*{!g&`-u��SI�}M�[�����p	(��d:�wVds�C��%�s��QT;�>H�o������ �^�A���&%��{u5:�LD�)W��Q�K��i�1;���yV-w��&����|�j��J�%��fcM�A(�W/��A&!74��L���޿J�m��^�2�ͳhǢ�O~���{[�(��f�0�.k���ez������e�+�Q��
���Ϫ8���+Ø�G�MNn�Cdyo "�-o�b�ܰuI���u��"L	>s�pI��R6�6��!T-�r'��G�(��ZQ�%3	�vi�li�~|���/v����~I.�*<�r6X�+�s���,Y�v�cȘj%�7g�*"��CG�#��(����@����-�jq�X�ޛң���-���ȷ�.%6���n'P����я~�$�,yM�}�X@� z�s��k?�-C&{ �^QÚb����`wn�|�QN��o߉�u�$�T5�IY"�Q���Mc�}o�W[�`�?��ސm%����h�-�]��hdEt��~K�$��vx��+֎�w+�ް��4��tJ�+��Str���t�F�y�q���C#6rT�@�J�ş$��mΣ�6��>�L�S�D��Q@��9�U�$@�-�v�cJC,*u���fۧg3
�(��;�.Ń>��z���$�x�gW���[9Ky��1f��o�{���b~����;��%	��X=���Ka<N��D�.h��#���y�ļ����^�I���g�ׅ��*�@�_äg�I��`D��k'OZT	�@�t�rSaSX�;ė�<@���$g�"����C?~�5&��ڣ��V<%��e+��̳.��P#xY��F��(�_�˰�uBFi��j6B�?�6��'�?@
�����91���Q?(_��x^�S�I��:��b%_����;�6Xٲ_I�z�֢���~�w7�����r���~��5�K����}$*$��>�D�ǽ6z&7� ݙ���(e�~�b�M�)�����?��Xi��-��R����	�ݱ�5K5��*=�~��DdCV����1�9�a�f_�[
���4醗}΋d������h��,�Ơ5�"鍻'��X��������.�DG'R["�aҰ]���P�JF�^�Z�׆�З6��5�jrW`%�#h͒m2w6;��+0��<�	Ѵ�k��|�<9>��H#�hi�ٻ�@�{9e#���z��%T�����4K"��hn6���#���t�� ���ӓz!qPNy>z�'Ⴤ�VR�}6�!s����j,;�Xa�wZ2"eqH�R�SJ���Go�	}͉n�������))h{����k2���Ȱ��.{�'�峨��j����C�ى�r�o.G\��I�8��,�^���	I�o�?>e��ڹ_g�}3�ew�����p}=��i�w=�XJA}�iK���=!]�
��6TO����e��e���p_�yz��?���p��� l�m��N��|ο%���3��U�����Z�n3F/�Qy٫�.a��Uki=�+Ccp����	�*D���	T���R����	�I�F>[��OF�����:S� �#	IRj~��f�Hn���UAm�G�r֜�clT��Ɣ���7U$�sא�l���ܾ�r�Sk�$���� ���M;`�N����J���%�w!H��'}��(-��L �f�yG���}UTR��Y��r�h�������C]��V��)bA��
Ηy��Do��(�a5:�_牤Ə�|����L{�c�z���h B��Jv`�E��Õwv�(O8!��6��S�>���0�F��T�P%�w����>�TH���.��*_�����}�����fZ��Y몬۴i=��y�$�-����� e%%W�{/��Mw�N�������������$����6��K��"��%�U�TD[�M�~_�QIΫ�(,��m�冱����T*���ŵBq�A+�%ǑZ�g�sF�v��"������h�_�X@(���[�vj�|y���uH'}��E��{-�zv��]�q� �������_ח�4گ,�1�����@�{v��K���D ���/�Y����A������x�l�oF�����3lE1G"�t��C���%�/�k�Õ] Xכ�'p��?�忤����/|�yڃ.�8�lĨ6��).�#!�p)&-�`<�cS�&h��r�*�3m�ʵ������D��WD�1:��`����[[�̟=��-��Q�)�p�����Kbrq�!F��>�m��(>|?!%'��B��(��b����>7v$�B�3Yu�����Ž�ǘ��F�n�U�Q:Z�{��fM���6���W�y�0���u���{���ұ#�������{��w��B�Irj���Ht�Q,]�x��AE��9����?d̈́�h��s�@S$\i���P����C�g�Y���K��~�=;-y��u1��^�~{
�2D@���4{\�|��x��Nl���3�u�:Z������"M�h������̷Qև8V���C�ҥ�3�����N8�{�L��2�G���*p}#��S��|cmٕ�oS`O�1��Q��l�6�R��A,-�
�:��{����+'�!��~�3�4�W��/bf�*( ��Ջ���$��V��[O�i��Z<b�*B���r��6�᥆�+��7Û,I�cbb�oI��߈l� ����g��m'^FO���oty����ˍ5i�s��$7�3��JFX�l!�쪹&�A-��-�p_��:�y�d��hE/�V�f��VCx�����2����4	ȫKƸ�9aUD�U�mRi;|��Iji��}���o�XaoINq����'t�*�	!��I���	2��Y(��U�w�3^��=n��y���;�X�GW��i�?��֦�B��z�J�>��9@z�~�y�����׿���s��N%8TZpLhrS�n�7ם~��7w^�Jbnf+��f��f��˥5���"�qk���"md�(�VKeнф5/ԗ:?���G��M H�\׷�O{�B��o'6v�ǢCVZō1�#�.�O<l�8�9������
�'���wD�O�T����m�G������#�XD��m/���垆�Ӎ�����Ƞ�~d�	!�^��}>D��K����m�Qq�1�Į��K�6���AD�Y��}��'v�m�'˝�/SE��M�Hi��S���!���{'{�L��7��r/����r��7���׫����#�	��0s%jD�O'��1\)�Vfj��&��9� ?�o�/�wS�c����g&B_����&�;J�^������|
���G����ή�>XS����g.��2���|�GJH/�e��CJY#ğ3&y���Y�IzR�������1�ػ#���E-���a6#�,�拾�0zU�0�� 3���X~��s��O�2�I�� �!�O�|n@̢�����Ɂ��?�=�����r�p���+��H�U؂�-&��!l�.�j	�o��H��~cƟ1�'�i2�-T&d4�4ӷ�Ѥ�R���ƭ=��������]��E@X��2Fn�V���VІ������i�Vv\�x)n�ζ���g}`���p��{�bחʶ������HA�35~�E���dD�]��R�#� .��aa&���Ɠ$��!�c�h]*"��EJ�[Z���ׄ�lK�57�݊3�Ņ_�hDXPII���{U7>=�ou��/�+�LLVjӉhԬE>�����R��x��\>,Ҭݨ���A7�����E����8̛�Re��1��\~�W�U�\�a�
��^o�ri(p�_ř(jݜ��/~]4>��;�BS�z���(�I���W��S=Z'�r�kQd�uhE�l�M��j��>�Q�&|�_����l��,�s����"��v/8�no��I�E�W[�]�Mq�˄*0���v��v���eһ�}K!�we��Q�I3�E�1�W��%D���/5S<���k�o�H��#zi�(�Jʎ.��u�'�W�/@�6�jq!-93����������G��Gn��D̘�6rE*Wtj#5�`d�OE���P�/�� �����	U(��BRv���Ф<�+�e$	w}϶�IUGHSO�K �ʐo &�Fal�0��{��d1n���/}����C�#3j�3B�q�Y�"�YhP���4p��ګ5���D�c`�훏T��eچ&k�]礜��wa!���^���4�+E]kj_�M�.$�8�☊j��ybm��4e�e��o�����c_v/|5�)��M5����~�]A�����M��r���}�M�ܹ�eA�>���Y�MB�{��!�8����sh�˕u��2�<I�/%W��P�^�:d�#� s�H�,8����)@��g���r�q����c��
-�A8?�#��5(�O�U~4B��p�i/�-�C��焤;�5o7Y(.��eXc�1vޟ��x��Pa��'��4��%�y�0��Q�����bFkS{����i�2Ϫ+˦��Ĩp�g ��])�t[���!������H�)��� Ԁ�yI��N���ǒ�Ui���u8R�X�����n}���S�DŤ�L3�f5��wX8��_{~�G'�0�s)��|�% b(PoJW1Fj�_8��=�d���0�Iu���ݚ�H��)��Ϝ��wP,76�]�?n��N^,<"#Q�7�4����+�岅J,j��nl����U&����$�=a��\%%)>�'�d�KG�{S��$���ʌ*�$[M_W��[0f�T��WC�P'�!]g��mi"����[H�~7b�0�����5q���}C�7s=�Ֆ�ڟy�Dն��]#�"3�""��p�7��b%
G�l���RM�6���{���Y�O�=>��u�9�+�1�����aAQfJ��aJ�����_ ZEF�ד��.!��K���/��r��O����U.�NqI��6�;�t;�땻��%c�0��>̝�2�2<Cݨ�G1���јS��C�<5�E�(Ig���;f�JLW��[4�+����#=�p�j^tۊ3�� ��D����/��`	v�W����;�Ş��x0)��4/��B�\�.�4��_�&@�-�p	�ػd4���m��u�C���5Dz��tŔ?T��g�[J���Z����[*��ؾkM+.}���_���$��[̆m�|~�H�(�B��{Thvx/��IQ�r�~��[[��-q��n:�$�N�Q7���6�� i�3�#��fȜD�S<��Νy)�:�<&��M���s���zgtV�V�2������U3G��cJ}�������b�fiB.�w�����_5��O�`* �!D��j%�4��1$�3��0#ѝ������*os���e�;��a$��6AԊ�:��w�bB�W��zlj����0tF�4�J��(V~k��-��T�_�]�'�ͦ��G�-OfIeDT���\L��k[)�����^~��.g>L��Q�ةaˌ�g)M6����\%dnH�9В��e�I���G!��	��(� ���Ou�{���l_��Z�_�S!C@��u����:�Ϲ>�r�
��-���O*)��.�ֽIO�i�p�q�$��˾���,�XsZx�Г"L|E�������à��y7��'o*�5s�Sf�V/�Fy�9q�t3��?��	�%�?}	�=�����z �����������gR᫅��eq���͍|/VĠy�:�3/ �cz>P��_�p_v-�L����|��o����Y6,-��&j�8+ve��B�i��#q�@�i��]?{ �a�[���e~E �u�(RW9I�Wʤa.�Ĉ�:O1�li$��&��(a���J�����ٖ�	m\�$��<$@f	Οm[&�;b�换j����B�/���ET����z��pB�|Y��� ���X�l��k����'��[�H�ou�>�,�ON���'�8,[֐��Dg�V6D4h����V�1�\K��q��g'坮����W��'�|\����|X�	o���j6V0ii��Bk�������Mc:�z�%jKm���2U�tt�%����3��[up7~����(�Т!�QY3Z@�S<C���;��.�\�s+ծ"��[�)m�:V͛#|˕Z�ˈ�D�@>a���n<���੧jv���-���O6nS+�#ф�׽ ���?���g�0��,|�.nc0V�)�~(��t�P����vpk:)��tIԞ;��C���yK��$�bI�%�������)����5���-"���g����9�`���v1}��'Sڅ�`�ؽAW���� �z?�.����o�� Q2<y��
���$��'QI�ŒL��w/�7�^���GsD=
-��p��o�3��>W��J�#�^5�s��A(��@PȆ�P���F}�ˏ��l%��v#����a� ��R �$����}�2��ccn�=��82����^mu��p(�w)Z\�;��ww+���Nq����;��������Z7Y'�I�ܙ={�3�K)A}N���?1��h)D���x��Ev��a�0��X3lΟ=߀�[�����Â6Zr%Ybv|�=v."os;6ːs��8.B�3~b،cT��n�τL6�H#�e�[���'«q#�|�NkSA�XE6��zl%=���b!3h"\C��{6�'�z�In$Z�%����zt�;��t��o߽8��y��*��䞷*!�X�ٱ�*�Koż'�����b���)�P�
ee!=[�1�8��-����z{{C(�^����M����ި�~��\�br�j�t�sN�-I��`�����e��x��ȓ/����OT9�z@D?w��|9f�}���km��p���L�,-����	��Q���]�N({�*^�����Ći��9l���v�P���6�n��m��Mz	�N���H�镅���#�-GV����
ѻ��1	����[�0V�� ͷ�]<�y�0S5���ɂ���?��0Lo�ݿ���,'�#��v�Z�������[��Yb���<�%gZ:��H9�bl0{k���K����j�iS�+��E1v�����]�q����L/Z9����4(�}���!O]�|��o�}�'�� jgԆO7�)Xک�l��i�?*{��9�6x���
��E�Ĺi!�r�-��??�nsB�.7�&�M�D�Fl2P>�p8��j;�V�Y�.YBkJp��.E�]���	ҏ�Ԡ�G�hUqGk�\yt�s�-�>v0f	�B��֖��ꆸy�u�.�r�,
;��:�$�}>F.��@� �c2Tc��S��Ni)9A���H��z_o(�:= r�|P؛?λ�jLpi�t�y�^NT���n7�T���M�K�e���M-�>P��9+6�P�?g���K��g'C��ٺ�F���o�$>2;r"W��W�k��	��݈`���`�L�y	�P�j?��T�9v�k�֏-\<�"��ڨ=L3_���y���[�!��SG${�"�ɯJ����v�#^5]��5���&D�U<����i�r;V`�s�
��{G���
����0����ބ��L�g����|�2Q�v�����}��_�炃=l��>Gw@��X᏶�C�{�݋p#��m��;fy0�>יw�&O\Rj:=�0ȷ�u�~ϱ��3�4�̕+{�t9�i'��)d�v�P���V���*��ظ�̔T������D�eP��F#7�]�>���Ǎ�Dԡ�ғӁ͘�����'}��2�r�2LG����j����1i�V�?"ѫ ���g^+��{3S�x�M:�S�ܡ�c���n�Nݖuۏ�(*cy�+:9h��{�d:��Yh�@�Z�f�Ew�$�^L�tԜ]�XX0h]���SL`mOB��Cr*#�hbӏ�-�w۾���nQ^�f���J�{1>+8��T��ZZ� ��Xs��c�{f����X��7�9U�cC����Z��Z��4�URq��eS!]4Z�y�eC|��R��� `�%�Ƹl��^Qg�m9����T��	&<�&��[�o��`���DfL�;MK>��n���g������V�bv�y������P;S�]�jED�p�z�&7�_X�6P�1�;U"4�[&-G���Ӯ㺰scN��{�YV�Hj�FP�;�+76��kw~C�^�ɍ�V3��p^� ͕3�?����i�O-���Wh]F~��[�@�<��^�zG3?����Z0#Fn�ܮE��<EJ�V2�bs<Q.���rV��f3�"�L���h��1C��)�oo�{�3:A-��z|��JutR�cpd9��7T������]�ϫČp[�`�Z�_޴�;��x�wϯ�=�WV��r��L�1t�Rg��3��	xd����^�\�E�CH"K�z��=Ҋ�DHI�����d3>Xә�PѨμ�yf�_�16~#F=V��/P��0�Y��Rjؑ��d�ӳm���y��ˤ����O��C��O�O�c%�3�o��iz�k/r؈x��%���SY��v��̔=��K���o���O8j�FN���fi�Rᩂ!6x�R�us��\��l����w�\d�4����UT[׭3s~҇n�ŗ\|�?�E�,9w��/�C��h.�����A����e�fb���$F��֌_�Ɋ�|41�+%�����::o	�K�����jB��_&)j@m�e�v\���x��_�@������0�y���g �J�b�lٙ�Qb��e|�bTО5���J�H�g������0�x�w�D��<?m�N�yЉ��ӄ0l����F�����1��5���=�@u'a��(.�*�x�6���_)q��͛�J��j���[���4pbBZ�����G� ���d���f�v���dN��\}�("b����Dq�4�`��7C)2H��Pغ�����'ע�ƕm�\�c�;p�%*S���?�:އ���ο�ij�㘈�������Dӻ�����`�Av^U�����y�Q�3���"P�k9�^vG��@37���E � |ئ��v<J�e!�F\�W�2  ���	P���h�U�u\]�v,d� 9����j�3�|����6��/w݆GK�������R���3�#(|W�6l�]�#Dm�C����L.&��>�q*�?� 't�}VRB1v�oɓQrѻ��>cyz�.�v�^Ptu2�F����~�����h�G����~�����L�^M��F���F)��8�? ����ظ�災#,��A|<П(���PV1@Jf����? ��@���ʘ�?���%6��]��48�������0���$�I9��)����vﲇ<Nd�C@�0`6��$&��y�[FQ�f�����c%;���ֈ���@�Q��a�=2O�k����%��N��OҠ�~f��%`U����w�i�_����{+�j嬎������܊CC"��'62�\Lv
�iSF�U<4q,}�?��'��B�`�Զ�ZO�/'?�@���j����hh�v��rh2<���N�e�z0ꓒ�nTn��s��~��G�t(k4��)S�R]����t?q<���o#U�b1I}u���u2��87��8`��1���S����+�,zv��`SZ�5����2��c	��B/d`4
��퐷�/^�H�0
�7��[�k��,Ab�`&��C�с�i	�=}$��n^���d�~��B��������*�����^���	4P�fI�D��}B����"j�Q�,�1�5�"b3�,���Ql��/P\4D"7ȼ��OT�������uǄ���I:�-���X.4t��L�7�*�g�j�Cq��f`A���(���@����*]+�����D2�O� ��$�a�ָ�R��@�"��#P���b�d� ��I�:�ݮG��ɱ��\;�ܹ�\_/��V��x�6ٕ��1Y�x�?��g�֜%BtF,�g"u��_�8g��q�(j��u��Qjd��-u���6��Z�R�#Ip!��(jE�ǃE
S��p�E�m�vb�\E�!� E6L.�����`��_�4���d��E/�Q��.�,�H�4�n��!&�|Swsc�yV����֎��k�&t��hi1dT(<;$zL���j�ͧoa���]��Mg==�����~V�M�W��"/�m��
V9��1�	w���4��9EP��C���ÑaC������k���a���%b���Z�
����������,�!��EaJ�_+���7?Z�{�S,>�}�^a�k�80��ml����O#�b�⿏��p���JI���o�@H�YHrr�_[��J�	#�����$�=�޿�)���>���gP�tЂ)N�����͟����l�������Et���� bӵ�mp$T9��{��)U�X�ʮ�`��g;�L�VA�Ҫ�Z�!	�Ղr���V����`1:�p"!n�
O1�aYmu&��f|HW)	2�d67��V�]`�U�Q�A��ڊG3!! ,Z���V���G��Ǯ�'j�����m�ڑ/=9;/���V���R�瞯8\Wk�P���>\.1k��Ng��f��a_W�J𳮢�p��Б�	���`��/Ɍ�\�&X�L(fA���%�����WNc&H�tC���i��!2���Z��r�Z��Y��=�l��.�\�+��-��$ґ��6�_��������b�R�;ʾ�^'������*b�#~��9��`����g}���V���HF9.d�����4}��[mgqtt�Q��?�9��ɼ/(赵����j���.��ʌ_�mİrZI�4�>��;����<_���@E[n�ڶc�m�
ϳ�f`��p�F��~�3[]�=m��[�d�"1c�;�t��l�����c0���������^����/Om;%]LC�j,�)O�����z����Ԣ�#m+�<}n�]e�ބLr@��Pf?��l�U|�<��1����P7�}c)��O���C�5ttI�na	�.����Yr3et5i9�o����'=:Nb�����s�3���'0��^F�^D�J&�E�{��K�6���[�OV�\�������P�Hez!��*Q��'�\���P_k����ls�o/Pb��͎j9�E�S��w�Ck���=����٣�C �iy��f	`�pP�p4FJ����lU�������7�g�r��L?��2g���������p��*)��R�)fAV��8��Fm���ݍę�t�ޚ���!�'rc��8�y�k��Yw`o�[8LC�)N�[���� �.j�]h��)�\���'p?�`��A����B�%y$�����g�����cT3ɒ��*��d�Òk�ˍ�1U��xl^�b��"M�r�Z���z)S];�$���}|��1�%��GY�XE*TH�I�I�z��N�w��I,y<�6�c�j��W�b� �*�x!�C0ʦ<��$�f�3�������z�xVC!��rЈ��0����$�;��͛$�50�ǋ6u	6��"K�l�梍 Z��f�^hF���\�{�݇���J�
W$�p�Fܿ�j�3�9�O�v
<h��5;�^l6�jG=�#�đ����~F�R�]�
���?�͓�(��w�yL(NY��{H�b0l�2�!�!��
Ж�]YAr�ǒ��(vG�s����}'���/Ex}�r�HTU���q^�{��[�"c���'�?P��;f�/�SY�_�����лv�t`�j�4ج9����+U%�,vȀwrd��Z
�~���h�H�>e+�� 7�t�h$�.!73�}����ľ�"��q�xí#1]�������Y���u�������۴j�C�!�~�������屇���r!�9�7YV2��p�M�T��/�"��yն��8�Efn�>E���2�1n��� �9Z��?��v��U������?�Yv����Ax��G�x?��.�6g�21,�bi�e�N��B��T��:٬���R%F*���9˝՘�G�d'A��dH,���dS�c�)�N��N�Jݮ�����B��?���6S�6R1�"t#I*u�<�a;5�,=�h��Ѝ���
>!u�z�Hȣ�2T��ڊ�p����]�\�}��\*���jSܴ��� բ��Jv�54�(��ڔ3�Z{03���8��	�~���#���N��V_��r�ӂv�� (@=�������n�{�a�|�$��t"8c��3"Dָ�-{8*��u�<�/2�(B0d	z+�y��Cn11��9�G���uؤ�f�Mˊq󐺀���о��L>�#u~g�5��'����m���:4��G��m0Y��k�_�_���<O���j��ck:� �9�fΝ ����]�!���0�~�l��u��m�&�
'F		hT���?=l�J�O	4p1D5�g�^�M,��m����łK9(����G�*X�!r���Z�zަ�c3X� px�� M���������G6���t�~/�Ux�빗�D�õ_<��c���}��*�f���o�����V�!d�:k���#=��b���⬽d��}qwG�?��q���z�=7�\s���pa>���yic��2���}o��k]����<M���E^G�$���l$_hp�?�äa!�x������`�M�,hm�=�G?\�	���|3{��A���i�#�0î�����q��Q)R1��HG�	F�g�k�]�oÚkٳ!J�F|LF2��l�Y����f���K�)?��v��	M�1V�;��7��XhYo�mP=�i�۬=hXC���$`
�(���	��~.0e�2S1h������";�Q_-�	�4T��}��b�\[$R0��H)�.kB��V�j�3�jeU�b��T�ɍ;��Pg�4mC�"�_��x=o��:k�"D(ɶ,/���Zѕ8JY�4W��\���� �6�����y��v*�����L�
 �r�k�������?�:Q�mL��w�R���HH�\��K�]��1o5&%[����D���~&V�������h�f��΃�i�йSn˄��g����}�e6�Y���ˁ����l���k��0�q�d�ď�:ÿ�t<Xz`螏�i���U'K�~�����ss���R�Q0�,�8�d�FҦ�����gw�Z}��Ai�٢SkQy6`��̻�8�ٻ&E$ɱ�[�q�V�!��q�� 4\�f�v+�@]���_�*�;��b��&�3I�rw�^8%��r*{��it9�o��0�����-m[M���w;�?g�Kψ���6B��BUZ��bd�	H��yc�s��*�?�.�}.�_^bT!��
�2���:^��s�Bl�r�� ¢>�\f�]�k���,���Y�&E5r�"������1��b��b��P���z\=�ծ>鳸�X���Uh]��f� ��qxx�b D�i�%�elDA�[��!�����!��i�|¤e�s�4f��XD\<^:	چL�B7�bd��֦m(H��ܙ���n�v����������vi��o��Pa/b�'�zI�s�B'w~.���t�o�,)/M!>���pIUS�יnv/3O�S4x��$����	I�ts��g�;o99]�*����۩��uIOCH��m�o�8rW3��-/N��D�L�~7��������l|S�ũ
s��]�7L���! � k���� ֵ����ID I���g�Q9�P��˿7X�;`�;G�{���O3�L�_��џ5��%���P=�[�rq�;��l�<OĜ�t!�Ћf��ٲ�S=�|5��qcA�Z`�KXD:í�1F0>T%���4똯�6�8�7��P�2M�����.FT�y|�����`3A�]M��KpX6b�6tC���u�dH���;K��9��������(x���M�����B"x=��I�Pl�;p��\ �L~�X���^�KΘŭ�%]��1g=�緍4r��rjѝ���g��9����E�GZ햁���L�� Ka!��Z��p:��ߍb)��������DG8���fg:˦"�>7��k���r�P���K	8f��{8\�^S���f�W�,�x�K˭P���H	�@5��9[q�]��%"��E�'w�V�X�o��D[w�nҨ��h�ݹ�LdzC�����Oj��|;�X���A�c��Dm�e�[�|�j�$�TCE�4�� �c�&�f�L�@��i]^G�{�C
�뿸�W<_J�#�dK�g�5/g��/b�&���VP* yC��;�l�HA`��S@1=�ՆL�e�gc7��v>��`{N[�a����jX��M�{�+�2�8�dg���-Q���)_�����W�zb�e��,�����:�r^�5���;�
C�?��ϰ$���4eQ'K���c�_�*��K�	�G!
�����ô��P	g�S�j������
�A���5E��B��;�L�7fH>1��؍�%O����˰���zSPg���&���ET/���p��E#�u�N����Q�&&P�I��)�O1^����V|䳡�e��muq�Уq��R�0��ʰ��+��ҥ�)`�]Ğj�bO���f�6�N~�f�u�`��ui�w�A�����A��m�6�CH@R:O|��_�Kk(M�k�ά�zRv!��pd��~`�~Sj�'C���Mq��Yj|�<��	��5��9 �m^Q\�LbwvGm�}m"�,_V�`��~�9�����rA���P���Y!HqM�L�.��b�g�j�P�:��L���NsV���:�R�}�Ψ�fe~n_����X��̣�z2����@s���	��k�N+��y�����M*(Z���tN��m�?��y�~1fd0H�^���^�Ikm9��1�=���1��g]��%��j�-�SY���ę0��,{��1W�3�C��
|E��s`����9=��~5��&����T��)�����v�L�r8�MB
�U��#�~���."�.��2��4����G�><�A'��p�����DC+R6�$p� i�~).���Y�'K��H�'V��v: �>�����u��@pr�.�T����&�Ўg�nA�qs}���u�,2��q�1it
Պ�ȥ�2�/jcq��hy�$~��9���@�G�J���K�������e��a��	8J!s���n����H�4���q���N��֑Y���y ����W�z	��n�W�l�������L���|GFU��{(�:P�I�]I�+z���c9�^�;h����|k*fx���6��r�0��Qb���B�;s>��������t��C�lE�P����UIZʣ^����#G���C�g��e���:��vb��a&��7�o�"�G�,,c��;���T0OZ������G[���۸�x�}Ӡ��g'TCD#D8�����9�l��/7�+�,'൚�Cy�r}xpi|e+I�_���MC��v�X<3cH*�;XA^̎�j���gr��D����s��L�鄗��D���k���C��~�97�qbN�W?DĒS67��5�w� ��0�uy!4T�/��b���� ����'kw"ˮw�����g�KF�.�E:áԹ�|��R����y0�T�ώ��4{y܁��zk�8<��󚸑�;"�}�a��U7ΜDLmD�]֟� b6�"'�W�+i�t���:��V�w��V���f��q�S���׺�O�"��6��;���:go�,���V�+��t#��~*����?���\�<n*MkE�	�{�k��d����vޗ׫���˵���q�@�W~Hu��1��)�hrR��VV �:3�e���Z�j�lvŧ�s��#�%o���U��}���S����+�N���Kt�)�?z�0��?�M��v�j���_���y~$����o�߂�}W�~�Q���N强�� �cy!��u�"m6�:�ԟ������`�4*2mD��3+��lo�qa�f��~��(�[��/k{��|a�R��y�c��"�
�rCw밫��Rh�d-�Ѧ����ve�h���~sb�l6�/�#,foÓ���<x���36��+��V��l���ҦbY�*�Z�>�R��!~MC����g�ԙ�uC5;V5h���𨿛���4u�ӽĄxLC?��4����g���c�rn��5����ݬ�]�7Ý!.��(J���T�vD�#�8�2�ݢW�,W�H!�|X��]�x?I).��������m����ڞ����J\�@;�_cT_��C��F��k��T�Bi��_	��wMX?�h�9��݁0)@��{�<vj?k�!|�4�IM��!�hȏ$�tB'�u�+X;
�(ӽ�����]��ܷ;!�2�l���6B�MO�L�P�ʬ�}�V9��g��r~:�S��PN��z��9m$�L��u���W��"V�D�w�:�����T���
�Bk/�L�ґ�ty�=�D�rBa�'��N��Z�j����J�C�d�?jH֜e{8Rv/�'V�U�A
�O{F��e�;Ĕyx>>x@!��ʁ��|Q�hO�� $F䟓
��]�t���IE�f�:�F���hr*�,qʑ{)O~�9�#O"z	X��Z��*�`݋Ta7�z+�͗��g{��җ�؋��КV!-��ҁp's��|���������C%Ae��wA�=�Bo:�z�Ɲ�}��K���b��^T�4���ٻzں��w�P6V���\��]�ñx)���;<blȵ><��<I�J���5-9;F��BC��o��:��7�uD�ۃ��x�D�5[�}�O�8�͗�E:v���\����a��3H;�|�rwU����-����C��M�Q�tKa���XM"��I���1�Wk�$Cۗ;��v�w56H˛yjۇn�}s8�Ϗ0����v����fw��z�N�zh�� 	X��x�M����*�̓�+T���(\c9w4�u/���dˏ0�P��'��p໌-���Fo�"���J��ց�s�A�s��}� ��-{��� b?���|�m "�1�A�}���U[ ��@�J�s�t���@�����3�Ƣ�D�B���r�2��l�P�"����6�2�p�'(�� -�rYK��r�y�ԑ&��j*ܕ6�Wo�]��6�@�����"c����óEp���>ވ��_�����9�X�4?�äg�GAA졁��&��jQ?$��1�D����ו�9�]؇�WN�I0�{{,d�ؘ�/�x���V���ը��7w?`Q|�@�m<�p�,�nOX�%�s=��b�"�aY����B�KO\%q ��oqU>��+����d���X������Z�v�H`�-��):�3����,Z�Er�r�$);]Rn���4��3�������u�tF�uwJ+�i�q�mD�jܯ��_�����NQ��&.C��h����p���O��%����˵��U�E2���VOs������}���N�2d3�����A����/|�.��y����N|;�+�ȳ�Z��!R���/��E����JaN����x�fg&��cK����ܛ<��.��tƪ=ļ������S�M�b��Qs>X�|��T�`a�_��k���7�����1X�����{)�1����h0#���f#�����]>���L��Ͳ��(����^w���7Oy�~�Fd�i����x/-� 6�8e``R�#<��-{ܡC}j����E8�  QX�+% u4��徵��� Ş��Fy�ss���8��q�����^YO d�Ӂ6WQ�xP�.�]~A�v��N;.
��~�m�y�iک|�v�rE�L$�Uv8B.�� Jn*�c�g��V��<�	o���%כ��wOȏbh�ǹ�F.jc�ݻ���;V��g�;�������]�_�J����GF���c�g[H��D��M��";I:1]7Mu�L�s� $bFZv[�����+`��d(������;-�S�"��@�I�QƖG�#ʋ1J�`!�T��Ґ�˒�-�˓@u���$��L���7�E��iU�f������*=�e޽_���Ȼ�\��@!���I6b�2���f5�8G�� 'I�p�1i��C�%Ռ��s�������v"��,և�D?�D�R��;��a�$��@��� 8�/���T�c'9w
����p1K(��j�ʅC�"�M�j��o��i����s���m%A���1�Q)��9��$���L]��dX��3)�������4t�BO?���[M��я�����S��m�;c��!-�MH\S�&��`�φ1���7���jh�o���Y�˹����G��<����^W$�AQ������S-zF���.�w�ԖG�a������,Lc�4��S2��gF3��WyT��J9��;���&T�6���� �c�`��;�03��k�����ړ��*��a�7�s�Į�|�wc��J�t}������ʈL�x5z1�_I�v�������SI�1+�o9�Jb�;*�l��T�9j�Z\wr�$9��v��u&��գ�t9�K	�;�; �c��`.�H���:L|� ��`:�Z��<���7hhRc��\�5�^�
���(Y����X�d ��>�����(|U�RD���ɬ\��)�ޗ���z�b��X��1C�p�B��x��ĭk(��<�����<63$��_��D2zTy
J]�[��^�)���ZUؖM�x1���#=�H	J��9�XD6���f͓!�s�m�#����a�G)�����14����o2��-{�i�acVc��}��	��X��Ea�a
��&�XNR=#S�o�[>�*��amxg��//���^>8D��~5µ.G��1u���t�����j�hj��#���M�X�[꛱HFnn0g���P�:�a��0��7z���X!݁-?��%���'ȷ�|,p�+��lhz��8�+̥���oP7�=[���+_F�2����8l��l4�Ud�ٓ��~�-�1������aq4oq�!oEm���_���I�(�/1��⨛�0�	�G�7���Dv4N��YL(�v�9��4!_�� ������`y4�/%c���r͇hR
��pDT찪)��k�e����4���>M�#��`v���0fh�Z�&��l�)�0��qp2A��X�#��u�k:/��Ze�Sa�9��;�m��������~�>�杋����p�$(HsX=Ey�����%�@C�
b���̖_[�B[7����'>(}0J�t���l���0̄�"�й�6D䩔m�F�j4Β��HvuZ������I+�4�7�^]��A�'##5�7O�M�T]_�d3��6����#8�h�Lou�NE(O��Ɨ�0M���3W�S�,��C#=C}5�ȇg�8��R��9�rC?���KE�V���2����w.�>3�g���#�X�E~jnJ��r�|��.e����b��n��_4�<Y%��۵���\a:�e����؎��_�M�Ϟ#��o,���G�z�(�� r���	��
������?���
,���@VZX~[����T��=�;�kl5^A����.�0����vR���z��:���,�Hx����']̜�oyK/e6�	Ke(�:҃#�i�ҲZr&�d52Y�7%����[ǽ�N��_�-H���!OH�����x����C=4
^�\��UN��q\Q�9�9�iJqG
�M�_s�=�>�^���_�z(n���d=\�0���1�Q8�쀢�f�A(�aLU��,L���<H��ۖ@�+��P��J��� >��BAr�VhL���Q$BCk��c���XD���yA}�î���oݥ����i 1	�����`p��/W�LH�a�vϟ`�}UoS�4N�-�å�>���W�ݴ���H�B�=���"�Zr��G���y�&+��q����m�GylG=����%J,����fG�v����>�&O�_X�D̈́�eS��8]/���0�tSk4u^-`���&	�\G��Fہ:�b򨡘@�>8P����g��"4'��U4Q�AO�CR1���>I�|�_T�w����Km�*3��GI6�0\՗�Un�����ٔhՎi���y|?]ws�6K�|���k?.]�g��0rع	���'����z��osq��bl!��������_P��K�r���s�x�N�o�r�݂I��N�<l��S.�fΣ�܅�S�knWI��op���&�A��{ԁo����s��#=;%�:���C�<��6�h�b+}�Jz���
Kо�Z�V`��10���>�w����
;���$�s+�:����i|G&�W��V��D��}?-;!FW0m�|SC���Y|�Y�n���8"���f7��/'�^� ���ص�P�mnME�}P��XWK����\�ʄ�oj(EUc����m83��m��ah�m�������@�`(K��L�L���x{��e{�b�ך(|�p�N���͈ɧ�B��~ȴ7���oS�s��{œ�̳�$YO]5��Ŗ-�[�Z�q�d��;���(�}���|^�@��q�A���@w6�9����#Ux@� ������������g����Y۲�̸���:c�UM��²yy����(�~հ�����e�^����
���èp�KLqk�n��j��w+�1������c��˅v�S�Skm�B�)�Ђ�#qf��i�55�ѵ�����&Y���U&�z|�7g�4��H�#�!}}<.S��v�h]��Hǖ���Wb]]� ��p��I�g�F�n�Gž\�oT�!�+�g��܍"_�%����2��țF�_,�1Gr�<�}��xk�X�K���~�r(�d�	�{Y�ho��G|fN���Z)�Ǧ�#de9�\��	;>���f`S����EL��U?�S��B�7��e��p��~w������SU,C�_�]v���jw�!��D���m�9X��i�@H�WH��~�����m|ʍd�~s�#������כN��><"/ �m�'��D�$���\� �?G��̙es5;�b�~3���|}���Q�l~'o��|�����08*)�Y�%��@�߷9��{ŉ�%V��ƴ��4����i%��;�y�N/���:�8.^����Q���f8�� 4d9���I����.{��5����
\v�y�������,M@�=]��f���hy�ԦպF5�����;����uH����I���:bQQ�9N�����ß��|�Zo����հ��k��וu>���ǟ�h%d]ٌ��5��v�	�u�i`�oU���|8�,���v��|ђ��\�4�LUA ��1z�r���!�g�Q�I�6��I<]�����[�.�9ʪ[�����M�f�yÕ��q"�Q(2�F�	�����˻2���·���+��bv�|���X�o��a&����x��k,g��d,#�K21��A,���w�Y�J�l�PP������JHj��-f�q���0?�6i�'Q0���
�%e���Y��f�~��w�c���;�!e��3@l$�r��׊H�ټ;�x8��(��6����Q���Z�Sl��X���ؑ���;�����!��Tj��]c[���4�+�ޒ��d��b�Kz^�ļ�=^�#���qh��n�Cm��c�r�E3�<s^�9&^	R���UKo(�1�D	�����z�b�dI�$��j�����>��E��@�"�4س��r�X��5˺�N���3��b�����n�v�1#c�^x����r��
�T�����OP_>^Y���T?M�EAt��{F���֧(�~�+�� ��Lp�V�!
)�t��/[Yo������(G��8O�1��Vd�1���	4��! ��w�tz�t��cqB��5�aZ*�jU drBi8JZ*<�f�QԮ���;{0zSQ�1q_�%S6��ׂ!'����ȥ�P�q��۾֡���?E�i_��x�Y3����e��u�_.�>�(B��D�&�X�Aj/��$������TTĊ�|�EM�W����/	��,%�'Y�T��?�i%�P�}C-�y�8��[ֵNW�+d����٤�#Y,ꑭ>���2Fd2c��YݟF|����L:*.��b ��3 ��i!��S0�!��'y�Y�*!�ɑ$Pk����,�]��������|�T���? J��NH��E�5��E��.�>��Ɓ����l�a��Oh�a ��ȕ]�ќ��>M� J#}dÁ�T�00XE&@'��L�V�X ��P������X���d��:�O$�4��&�0@|����r����x'u�ǿc�dM�yZ6�z���fZ1�CI@�R��=I-T#*�$3>��
�9(a!��	uZr	�ʨ˱Fd!� <=DQL���c��>/�Ke<�)�X��-�_9�Mit�a�PkSjjLh�)r�K�uW��
F��R�[��9�G�ɝ_ğp�)(����\������Nw"�����Qfrg��7d�y��:�S�nt�� �=�V�<]���b��x��2�-�)��Zp^��J)�D��<�8UT����H�+�p�"JC>�Uy���A�,���b��PX�f�D���:�h��ݎ%�S���eG��jUQ�5KŎ�KV� ��gv3�K>T1E4g��ZF�磙~gME��h�$&n",����֤�7��ݙ����3�yz?��'���g�)�X ���r��ꆪ���*.���琐L5��kƪ-��:l�b/%�l���#Ʒ�P�N�[�*ʏ��@��Z���h�-�x�)7� �"2����V�L��/P�~+7���a����i��Ԇ@�����4��JE��N�.��g�|r^��g��î[i��'J�s�<�p�~��*2O�F���~aΜ�g�Θt��@����jrs��j���F����8�,"� �?���-�&p�"444 `�B���\W�]�dB�=L����*È˔Ýd��!	G���)�����G�;8G��[�Nl�۞L�L<�m��$۶mۚض1�3�w��'�ԩT��;��׷����^)z�d7�Zt�M��K�7$8���\B��������WF�%N�DS� �W��gˉG��k�fz׷�#"��dz�d�`X�������wM�ݑ8C���v�6R��-�=Z�w�jڻC˄��!q��@҅2����5�a,e��f	���G�z�oˍ@��"�����#���Ju�A}�9>..�ޞ��'Z8A�Z��tx���G��<��d:[�/u+�nԉ=����Jiee�d�8x���_��$�P���0�mb�!y�9A!�/�S�t�
���
�^$M�r�a��00 B|�k177���H
�%nh*L�v���T��dtl����RmtrS!@X�б!�;" ȑ�bM�(.-M�׸'	��K�L�K}�Av0�$��G"'���UW���LA%��eg�{�`G��-�����u��BW������?�Ч�4xRcLW��w�[|cD����B��y�� ���a �T���D�A11�_�Ӑ`� BHJ&����,T�S����НVſGW�2����s�ϯ�0��:`�)��j���)��Z�Nz0(L0��7�熌."4���p?&�>�,���O�x@���O�C����as)I��7��Ȟ��`�K�qN],VM�!���N���DC۪ʈ��$(H{OJ|�+fۦ���o�����5����q�˙���W[wnM��It�Mny�r�U���AVS�"(�<+�ᜃ�t<�����]�xu��������锭���s�p�"nw�D@�nS��SL���i P�3��M%:p�\7TAE;��jR#���CRwx?-dp���Zz̏&0�4t��o�r6���}<O�j��
���7������}j�NM����'b �YDpz��eӝ�����#��I+���;Pv�'�e��󖢥�~���Dڵ��41M!+Ɋ�?���5�i>����J�@�1n�������s7�|A��O�A� �O�P�-�k]%r_�ȿ�}@�<��k�p�>����rk&�ҹ��ܸ=:愶y��9�QL�-�,���s�(a�J�#뽆2ಀS(?႔��9�"Y�h!5���$��E����h�y��6���H$�(P���s�2��y���Xn���c:�y&F}�)kJ+�r����-})۾�O�,��2I�JbP�\]��(j'�pJ�̂������e�P���w΁���,rU׭�rx���M�,��AO��$�
�X����A������z�;���8c�g��-w6�(��f2�+��עc�3ݞ<;2�J��c�����)�K�ժ^�S����|m4�y��	�������/jZ�%A�bnU��	nJ����Rڽ׺����ng�O��/-���o�N�]	�'���Jܓ�^M"MD���	�ь[E�I���<v`�o��f3ny�9���3/���Sc�BfM���1N���4����ު͇��{��5<=�5ng�;0��{��/ 8O��v���?r���r}�����AwȦ �)�����`���=�ʛ���'̝1��J;�������:yH�ߙ��r�s���,��؛��ճ�$�σ  ��'�_D��G��@TQ'\�ϊj5�V�8����?��e$R�7^2n񻽵�U����[3RK[cI������կ�<�.��������5�7g*{ktj*?��h6��S�#_���9�� ˡ��;��D��~�"��JW�G�����KR�Q�z��+E:[d��E������,��)��tٰ��ӏΆ�d�~�8Tf)��uxh��I�k�q��4֩?N�c6��^\Y�u��]$)���K@5d)m�X�C+#4�R��[`�T�����0���H��g�S�!����r�ѶORc�U�ժfG�RLm�����uآy��T���BqdP� 4b	Ԧ_1A�:��$9�燀��L�y�;o��[o�Ȱ_��r�a�^9	���NKq�&�0��$��NmT�����5=�����M��y��X���r�saJ�
k5yM%���d!��5���`�8Z�.3��ǄS���H�P��c1��݌H ��nM���0�ڽ_.����[��W VȞ5�?ʜ���/�#zp��"Ew��&�cE���'�PI��4����?6�n��
��a	�"Ǹ(���="���H�{-�C���B����)�YO�j�-��7$�B#�(Q,8HF8�D�F8�`��R��	υ� �#3���:�q5�$�j�ҽ��a��tx�n��{�<^���QJ�@kw�'X����p@�P�3=2Q�O(Ø�0$p����������Z.�6M;��k��o���#; ä�C�^�ls;K%d����x��l�y�-�Fu�
�寴-�T/k{G�U��«̅n�z��-��m���L&!�Hǭ!'(U��)bte�#��H`�g�	ոi�����N/��(H��grњ�A��X��"�B�� ry=j�I�互�}ۢ�?@k��u	QBw�[i�z�;?UDA��N��N�l�{~�9�k������:>Z�6��I��
���`p,��N�ǻ�+����rWv�1��O��(�������3Ո_�u�I0+M��~�+B������~�R�y=� a5<*t<��D#*�S���N�;�4^�����D���&'�3��rN'�B�m�@�v-��rPz���0�(r(w�Ǿ�E*��W���3&~�Ab�[i��V���ѿd�m��a�b�I�a�J�.�Pi�^������m� ��s�t6WC:�3�!�m^G��lx���.�J�[WO���0�ѥT`(�d�#�q�q|���R�� ﻞӾ�{B��z��f�q�yY�M'6'�«~!7�&��ϔ�tCȒm���k�E��ԕ��#�0Ps�W���bbx>�V=��=�n=����&Uz}���5�=tc壼�wC~}��Q�ߤ~7���>�4ːW�7W ��E� *������q6��)A��A*���]�RV��~�JA�C'�9ߞ���rșW��U;��*T�cԀ�b���Gĝǐ�����:�fWo�N�HK-y���MMd�q*�忞>���1����w�pq�[%̞���#�_�����2ZX�>\
�w�J�3O�����)F�ۡ�UT3���<��Rf����"p��RT�0�+Lǭ�3����od�P�i��Jwp��"ֻ�@��N79�ņ,e����~��)J������v�xY:�&�-AFP|��F0gR4��$�ȓP��?YL鸪��h��8���e-��7�h씵\&�j�:k�*>��l�T����C\���B#�F�!6ϩ0Jh>N3��6� �H��nO[��6Cڶ8�F�JL[>���;ο�h+�0D�g��`�����@^�3�͞s��**���_�h��=ϡ ��4M}�� �s���a��LE���DNZy/�A��+~t^*f�ʇ4��T��.�OˎY�������,��(�E�g[C���4i�hl.�M����5O�����I��8��PJEwx=�gz�k�@�UF}T��Y�Ш(�� ��r�U�bJ//~:M�^�*Uؓ>���r��FZD�}K����9wmT2RnK�Ȝǯ� �_�l����ƣ���/2.��!����
y�2�V\�m�	[�'{�� �v�*Zl�?�����oq�K�|S)YY�ۣ뛛�Ώg��؉"N�)\5�)���b��]��~�{��?6��\RbC����
2ѯܰr�������ch�U�b�+u��8>�ө�� ��e��y�7�k%���s���)
&�@gp�ٮf~ُ��׍��xf?�<���.$���O\���b���ܑ�����)����{�T���yhS���yݢ��[O�S�5"�<y����딁ɜ�.#��Va����֪��
f�`}\���#���	L_�hEhŵOZ:T�7n�'�F�]��S��ElO�B. ��JO8����8Ӻ��z�a�����Ew̓v��ِ��*�z���~Ҥ�޲!Ve(����q����.=2&���\�E)C��j~A�Wւ_u����N��g�W:|	Gr���%\�j�x��s>s��`H�����<Ʈ�6�X��Kz.�	.S���&��KwҪ��kk��<��u�t�����HLy�����YN��]�d�+qԅ�-�G)Ygۓ����q�X[����G4�Ap1���w��B��O$f�9�-6Z��Q����S���1GV!>�!~w�POĦ�����������+�|mp�f��/�@��)�*�'�����$����Ĉj5�ua�q��/�,�Y�����\l��:�/ PU�j��E|c�bHK������&����㙞��T�D�j�)*��Z��^���gO#�t�7A؛:
�|��F|Ԁ�Ä��C��@)F�n>�ڄ����>����t!��Qw����TԖug�����X����A\�I"�w�tx��D��]V���
�4�1߲��7��h�5kt�o1�@��i��^�����K�\�u9qq�;}eFզ���*�b�6ł�I�i̢(�Cre�`H���pjۜ �@��qe��Q�`i^3�!�V$wS���V���{U�y�� �Zv�<�Y��"h& ض��\��|�{}ɼ3�%���avP���P3H0�Sj�A:�Y�Ȗ�{;ׄ�gO-tO��Nv �ݡ{����_� LϏ-\��XGX�N�"}��t��t�
j�X#�!7�a��o�5J�+���]�۰��:!{}��ۿ��k��vٷZ�-�����>��y��y��w|-�b&.Ī�8�٨�"	�H����b �l$,�G�
>��7ՍF��m���Ȱm�h�_]�_��Pud8h@�~��~T�7�e]�dltHQi��2Z� a�lU�1�<UV9Ȁ�^^�c��wB}/��,�~D�.�$�Za7sR^��uםJ'�cӾ��5`@�:��[�����[�6�x�����|P�& �[W8A=�e�	zz�jX�*~��HJ�
�ozȱQG	�G�X�Q����H��}#�ဖx�ʸ��Z�P�u"
,z\���y�>����mx��\��o6����z4#��ޓ�*a4M�s�xr#���Ø�{yu�"���CL�(��˫��LE�We���ؖ����39�֖�3u�s�YWo��g�j8���P?���׶|�M��c-9���Q��f��e>�?-�#����93�}LNJ���4tT"�����%��x;��M���;lh%t��%b��s���\���=���;2��Î�ﰣ��=�(�	��7���Ǫ�!:���Qs���YY�Es)W�毷���k�
D0��� N�����hk�ʇc��ks�>�� �Xy����`����]�؈�KƗ	����Z����==.�h��`�H M۫h3NK&�O�hOP�X�T�ގ����jM�׍U8_� zA,8Z8˷���}�RA��c���,�s�}�oi���W��-��e|��d�cmפ��]X�i�w
�.�M������e���I�:r�=nx0�w��[���aA"�|_2���v���;Q��O1 MЈYp�?��zA�"T�/�Dbx0��F$**�"V#�D�=LI�I�3N�XC	��@D	yE&�����#�πC��[iy��L;QG��)a��F �v՗�(@�XV�0JI�)�uM ��FB� �E������lЪ����`X�ӗPJ�D[?(o�;:�3L�7���9�O�0
�]C�1���Ֆ=}�	��ӫ��^��R�{��L�t�؂�)�E��k�iH� Y�Ux�
F3$j��u9@Rk2���ޓ��G�%���,)�Ë�S����,���Kie�8��v��Ap�)X���f��d�0��@����N>	�<]?�``��B�ŉᴣ��ܓ{�2K^��m������q��謝B�����L܈�ⶆa�P��߁xo�n^��6��<^���K|���}�݁W?���3�:�TH"8߆h�J�Wy�Tw��[\�?�e��@�w�%]�Tdq��'�QG��i*��ǔ��A�8�QDR���C�n�n�@Cdy�vݸ�%$$�g�\�ʛ�P���<=3�	D<(e���/9���<�(V��}�D2����L��rL���������(��S��2�GX��p2�b�셇�E7�/r��c�Y�f��GI��!L[��o�k�)r��z>�:�/4Y�wuc1��mp(4g�"��W��r.�P��/�M�l�2D��ֿ��EE~�A�+Lc���7��4{��[j����U��84���17�������y���l�l+ڟ`�����
����)"��,���O'��ε�PRo�]��@/W���թ�����?�vq�����sf2�琣�ۄ�v ��@����,�~Y{)���)��C����g6�J�qY�	P�Ы���r����lo�2�ϛ��,Qt�tA{�6����`���彤|@���|��ha���!�AK��h:x��$��$�!q�G����U˙��Մ��2�	�3��f3�K�z`�#;P���dmփ��qڗ�f�����aQ]���c�:���S�k]^�졟��M��P����D�[�B
��b��VY?����a..��-���ׇl�A?�A����0l�A<��2�t�6�}v���3-M�-O�H���.H�ޏ��ʫ��L�'�`B����	�$H�/k�|�k��`�XdJ�VKgL׍
85�����"�Qp����n!zkVV
��j��PО��k/��غ�ۺ�oۺ�2��1&벦������AA�� #<�\�
�b���!� �Q^��yP�f�g�_� �lE6����5�N" �3�o`�E˯"�/§s[?�8�)O��2Dã;ER�Y���R�'��Ƕ��N�R4����Eט8�1�k�3T�'����=���ꀈ���ZZb�kRAX�V���~%���$Mml����`l^lDA��Ht��!���	��͎�0��a�_����+���L=�-m�*��pÙwE�������0>v"����-�U=� ���j�5�ga!�s��)�($�u�z�i��0�����ˡ>=�*}k,��:0��V��d�H?,ʳ�MZ��� ��Y�pUm��:27+V{��w�����.����@/��~�Z�@%�Aѻ KRc�cW�w�ͬh�:�l�Ze(���+x�E�<�&M�8Ɔ���gp�7��y���� �ث���i���3�?׀Wؚ^q�9<y�<M���,�k?���te�7i(�AԲ퀛D){fs�_!��t�+��W���g5��
�=� ocQ!��N�~E�8my:k�Q<>�8������^]�[U��HI��v�ޣ=!c��	k�*-��^���<�:-�KDhg��G�L�|X��R�YB�x��2�#1�L.��E�Oa:�]� B*ߪ���]���h1���U�S� �t�5�`©�:���mEl ��ɫ00{�J�Ʀ��8�)G½k�(y�?����lgr٢�j ��w6;��{�4�L����!iŦ�h��EB@e��x�粷�c�5����5�xY�ph���~�awN�Vy���F���6�H#s�)�!-��(�cւ�O&�eۃ�e�B󭨉�4n#%UUO��`��E�ā�3�u@ �1��p4�U��^S�!ihp���r��;������cҼ���/{v��$]�:�H5��p������Zt�&$힤u�φ�`k�����%��+g��)��v�-R^P�*�����K���;�g�F���<��h�v���[���f�|P�M$�Q����|��@(�0����6�m�>���{�q7��И8Q�Y
.�o���R ��h�Bĵ���st��|�Qb��?��ߘ�{�.hX�=�����(.���::��k�s����[�fE1z���^>�v9=��RQ��/���8g�|��t
���b��@�x�n�����9w�]LY��^�5�iw���*��,���m���q-�RVȖN�W
��3��C�<�/`f\�-C)��qwy�B��Seg��)��q&��Pd���3�S�Em^˚Z��a��8ˌT+z�ĵ�
�h�웠�fod�}�e%�MC��zXմ�����3���֢v#�x^��D�L'�ܼL�-M�n��e{��`he�d���W��'}�����)���V�廤�p-�cy�AZ�*�@�ig���r��y���ǟx�2p���zjq{�/B_�`^�G��!�����AF��a�+�VM����lbx{KRl;���K1+��.�8��6L2��o))ю!���z���Ao>;��\L�X.v�nF=`��"a��X�E���������]xї[ލ8��_sB�K�������Y��̵��U}����D�ƞq0oU���T*�,T��h���,K�z��0�Fw�x��򸾑�qލ2�G�G#��Z�u�r��M�Q�"ybuT[D���x}��5)��I��,vt`�s����'�}��H!�~�&�AƔ���,a`�r��k�1��O��4��.����i�E"]<`������ke�#�X����iZ�����ܠC�\�=j�g��g��.���{�JO�c%��~��%`hԾ7aL���ep�����y7(�
��`'�m�`g��=YF҃Z4(C!�+�g�����/���NC_�d�Y�X<q0��ԵY{����%�h�H�qɿ�K��d7������ś�x>�_p����6�%�qy��=��RQ���Л0�|%�������ƛ�}�/�-;�	E��P}���3ѕ�������u],�>���?GV��_�?�Q���B����n�\�z�%�Z{Z�=��v��^���;���"�W=�&p�\csR'Uy�װy��y[�<7�=tJ#�t���ɍ8��Yq�K�D�(:7�~g��JD��fپ'�,V��|qdG{���[y;Vc��Ʃ��}����U@�76=ӟ�g�#V!�dw�y�����D��kI`le8�u!a����������GZ��R��-��N�՛���"u3<3{�<��QT�Ѭ�.��0
��I^�K%����K+�I��O��� a}��U�1�-�G��E�l1'AW�ʪD8�<�όe�Z��i��,k%��5��=�&���cCќ3���Y�m����ug1�Kw�ԓ\n����#����m�ࡧߔ�A�� fo?	�o�`��>�-ZHru��D��ޫ��J]o�B�T�80|N5�?�	�7��Ej��|�-����&X�a�>�>��ML�@8�,���]�I��ke��K�ȡ�����Au5�4�U1}�Z�z�#;zpB;� ���0�����Kt35�l�����^͚��D�>w�
���3���v͹NсQ	��wF�P#�w)	�?=���o�%x��z����:oYh��6�֛�c
qE5��U�`���2��y��`s��}�E9�~' ]oo�
�֒o��/O����RrʛI|�tXRBҁ���Å	�vhx~L)��[���߾�G:{,�]�.$_�$5xk꜏�q�N���*b�3��I�O�j����R~W��N�E_����@��c�^�ZFϲmS:��5�*�2|.��W�@pL͂q�H�_ݞ�X�"՚����g�1��Yį��F�����ґ⤎X"�;ԗB9Nq��T:��ј�5�r6�J� ��mW�VΝ��V_~���a1� j�
�� Ӟ�G���D��d���<L��'��F^�K	�;s�a�%�  %�vc;�{y
A��a�,�-�K�tZ~bQ�H�"s]yu�Ԫ筂&7��ɻ
ѽ����"�/�f&P:T����]�I-�.��y�P"���t���B\n���#0Y�F3��Ct�϶�AD�{dM���"h&��48�Q�q��s�,b �3OOI_�NK�m�·T����z����mw�2c���	�;�%���s�9�Z $4�+Xg��D94�9�RM4(�Л_��?��3U~�x���J�밅����eb�4�dʀ����;�	�yD����U��(#7��[�(��f؛���
N���9�ԁz�?k��Eބ0U��]H12\�⣔��vf��X���K)�.:͏�7�ka_ӊ#>'G�a�Iǭ`�|n0y;oH��j��"��㎯��v,a���]��N�mc�}� �#W�.���
P���S*��ùD��ũ����rdQx�^�_)s�@��9��:�?�*y9���,�Y'囡��ņL+�ni��k?���O0��9�y�?�^�@q�b&9��4z|ϻ�GW|X����h�^_��7���r�k. �TJ����ke�af�y�̊���ti�,&1���<��Ac�����5��v��o�N�v�WkQ���u�m����*-�ɬUD�˝��`��款C����Q���[.�������rh�Lt�-��w�� 9��dTR�!��%A+�Cڗ]Vْ�B$�fށ��M��)�V+�ua���{��5>N#�Bqee�&��ZH��~Źa�П@��[���
�3�.��xe��;����wwo��)D����8B���{Z��N?:3�h�x3��pn�rC{�TZ
��Fy̍��RD�ϱ�6^�����
hX���P_�,V؝��'���Ʀ�����j$�3;�q���]bȊy]d�\Y��+���n��hq������-�E��c�Bͧd��飼�H�Ƅ&zo�� To��"�g�L,��X�)�Բ
h�gn`H�y��<����GR@։0���+�"î"��P��I
�X��܋�=��0����9%z���y�m���k5Н?�23RG�V`�9,�?�L2/U\����49`f+��ׂ[����tQm��:�J1�9⵪o�S��߲�:���b�AT���ɟ�%w;94�K�"�?EM��q�����4�����6tmx�Mt������2= `�� P�jX^ڈZ* 3k���TDd 5Ԯ��t�S��'v	�ei�|���������VNQ�n@�n���^��=���զ�Ǎ5o��ea�&G��!s���J|����{��)�F�8 (��,�/�?eWhl��ZE8/�v����I�r�}%]o>#((\�*#˪V&{\z��T���%N��Ö���ڱXp� kW|jI�\�0T!���R]���t3`��		C�y�����K�2�A���%7�[��	��ӫ6���;�&Ƴ�& �="(PZ+���\�-���5;nZl�#� ���ٯ2�:��A\9`��5�<�Rjꬻ'�Z+�o�������S>~�K�Pkפ�K���/���q���tހXk� +t�����BSE%�r�[�嵺�S��\��C|�K<�Q��E6�lGT���4N@�SJF.�?�5��<��|j�W#Б��sd�x��r7�)�To	�h��+�'U����ipf�oң:@k.�<��[���F�˙'g��J��{ ��a�\8)/��j�l���-��Kd44�]�	~�e}���gKf��.> >D�t��Wv-;�	�y����B��8����U{#6]����/"}\�f�}��hR��(�̚�w0ye�\�^K�o��-Nk�z�P��F��K'΅��dJ���|@`���V`�&[�
Rw7s��7r��vP��dĺ�Kwa�V��� F:[N���5(��2r��;���fhAa��#�~De�n�?���;
����fU��;@��>I��9�3c"?u��{J�w3rV��+m��)F�i�\�U�@`��MZ�$�l��2X[�-��E�V���⡁/q�ki2 �1�����P_<z\%��<[����
����v��!�h�t�ܐd���S܎`�$Svtkqp�L���e����&�4�1�|ֈ-�v3�db�71;����\ǒHp�zw�3(8�$��Аa���c�B_�w�A�$(���,��׶�hf���})r8�3���f�hu}�~�G7� �7[&^�04�ÆLZP�鄗�[+�Q�G��]?��"�}��u�0L���9�c�{gc�>���3�?�)0�(1u3�� �wsm�7��Z�wb()UA��VNsΈ]��tq�_�g(��j��{x��t�!�WY8�.��G;�����z��|9vo?�p��Fv88ӴFq(��oNNl�*^]��"��޿��nv��"��E��SSm5|"��ĦvT=bv�<���L�i��!1�E����(��]���r�nno�,�Q���g=|�fϧ�؏�U�5�\��0|A׷���YY� ���xVZ�!�@3��;� e�3�ص���Ъc��z�#gi|?O�x��^)�%!6�gO�G�"�n��V�gX��
u�.�v)W�7O�-}�΁ZA?9V����J��rfΩ���B�wqU�?n��F�5jp�it�"y
�fO|�m�R
�Խ�=��������8�Sӕ�0|�er��ዋ��H�u�iJ�X�I���5L-��c�d`�3�2e��^^S�2#�c #n)��"�|�xu��gz{;1�uZ��X��ҭ<_\���)g�D�����@��ո_�)>TA�|��`��L�i+��o�҅����8Xgc�K0��B���컷M�����]��Z��7��Ƙ/�����2$�{B>���ϔ�Бx��/�"���3r��?*�_��Z��e�Eř��� �G����*[�'T������_h�A=�h����������3s
�7�Ӷ�� �\�!4_F��J 	&(6)���K�Ǐ��ْ�Q(F�5᭼�si���g����c����۸�+�'ʗ��^�NpAs�Y�:��Z#E�2m`g3���z��	���P��dMbWCIP�2��Sd�HB���rFnlh�N��]'_��w�טh� ���ݸ�D�B�=�P����\D�E.���`q�2�跴��M�AM�Tp���5�������%�ʪ��C٥#br椊UB� ��a�7/��y9ό�c�zp@Pm�b�/���oT@�ș��55tj[e����%q1V�&�՜���(�����k�rl��}�VٟaAQY>���` �4щʹ��Qr�?���Q\N[¾�(V�� ��,:�o#.�-}bǦ,��,����w-�X��@�t|�E�Y+����]ʬ6�n�w�`={
���R� !��8�'{�����U2\�Bcf��x����������#Q�N �i'�?���ܪT$�	cM��#��h�7f��$8H�B6���\�.������ɒ׽iD���ϯ��Ӊ荃�V��@6d'��v*&��,%��6�9�U%3��*�J5��eȚ�x��[�z�gz;��(��#ܥP�b��C����7��?���q5o(ʹ_����-�V�_X�Q�p�}J������v@�?x����{|���˷wE�S���3S��b�U9�̓Y�P�^Ʀ�&�
�s��n��P�Ow�~1��g2��Z9����,��M�X؞ϚSz�<�Gu%��z��!OMG%r�O*�����;���tߤ����չ���Pu,�����nݡ��r���̈�����2�p(� hP�o��Z�6��r���\bcB���_W�g<��N�3w�ji���{t����Qt��GEv��aVI��1����v�6#�����Y��>�9����ڏP�?��z~{{���������3��������I��@?KL�kǸ3hlrÍe7���ԽM��N��ZY�f��(��l�x�5����.���y%1�G�n�H��J�����
M	��ʛ��&=������
+�+�����.ȓWEjtO��!;jo�i�VO�osC��ʺ�M�\w�?�^6�`Jw�q��J���!z�K>��w6C�XS�HG���ٰ��)�A�XJ�3g�`�������1)w��˒G���ʔ�6��Ė�G�]Q�k"�7,-��o!� p�v��Y�:z�Ae��𩈪��1�/��<��5>Pp�o����!��Υ$A	�L�)j�E[M�1�_\�덌��<�����=eZ�����qB�~^�;O�g���Uwp!J�o��&�k-�#.����r;���ɈtcK��lG�8Xq���5M�YK-���q��̙G�p<A�	��0�{ ��uEZ�/bŗ����*Mͤ22;�w	����k�S K�o�[� M#��� �B�W`f$�z�Q^݅�;95T|��:ŘX��i fZV�n���Ag<���PAiA�]=&��Ɵ�6M�n����Iz��7
RR���O5�ׇ[��$s1����k|����X��_s>FQl�{V9�o$��R�sW#�-Ʋec=��2:�1NT����RD���Ԙ��ٙ\UT1���&P5kX��b+W9��b/�-X9���!}�~}&�
���zMi�8���`����Ф��X\LS��eѸ~���n:�>eT�@� OQZ�
���@0s�?���[�A�괗QS���&~�nD��/��L>[�(��
��1�M|�6FVyA���ݔ��w��X�IO����Ӕ�l�Ϛ}��!����Z	�]�{3,�D �E�c;cn"��&�j���sa���`���?k�q�������@�y�Eg���F����Ќ�Ys��r��efm�h�̭t���<7�6������۔dQ�?:�]VP�W���B�i?������(�>-�p�p=#$�.��ry����j[W�Ī@�C���;>��t��/�(YNz�x���#����Q慄ւ�����\��	�֜��|ǣ�H
B��ɶ���8�O�6b�x�v�f�8���ŧ(3����T�1t��ߠ�fx�Jh�Z���%zc��m6Ӯ�R�C�c�tB��Jz|����������ٝ*7;>��S�īQ^t�Z���oN���,uΗ(ޮ�-�W,��6/<
]����?8��1h�j�L���O׀����,��}@��d�to�5����3=�0���}��i���DUbI�<>b�݇%?��O�"@_����X�;���I/Sݠ�}]y��h�d�x	�ͅ5m;5�����yϱ`�1YV���������|}e�#ۺ��_�D�3�+�mI��zh��˝A�5��Y��o� ��l����7�K�j�������J�.s�5�pQo�DeR��Bc���%����ޟ�����$��U�EM������� w �|'��ʀ�����)Z��N�h�jdi�c��]��χ xZO������:�]��U��J�=5anΐA�ͩ�aB�j���r�s��G)&��D*��2P�C�B��w`�
�Ӯ�2Vk���̆�D}�|��=��Fׯ?��Ա���`8�L���������fs(����33rM2<z)L(S�o���׽���+�w�D�7�<�����CZ�s7Q���)�+%|{��v����mS��,{����O�U��̗���,�z:_H�ꡉty�C��I��OQI)Kh!�:�PU�ʾ hS��֛�n~��%��q���U>D��^����z:�Z ��;}Q�}a1�n��G}튇7D~H�5Xh���x�C�����9��w�v�����.�|�%cr�]�]����>�A>��fD��J�'p�2����O��(�Op���ւ������J-�|SY�zyq��ύ�:�Vx��Y�o����5����6�K����>��{5z'�`p)�L��L����r�u)���R}:��h28��&��'=NJ���ݯ%$��Ba�)�#Ӎ����r!풪%�����K�*������ o+�U�q�0``dw��r�T�lھ�%c��<�]�R9���t��� �G]�R��V�6�+�X�j�nՑ׍����]�њ1�.��͞�p�~oN��y;��>��>�l�GLw�����	'.�ӓF������E|.�kQY�5����d��	�M�ھ�t�c�j��Qi��C�p���J��wO}Ԗ�_j��}��)�_�X͞^MШ����\����./�V�;k{�¾h�g��HDȫ0A��]t��U�2sl"!2䘪�1���
��:N����8|��j.k���'����s�Vw#5?9��u�t|����D'�C�⑺u�h�A(�%�c ;8��1]dTm��hp��e����^���5����9�H�7�wSf�$����@QZZ_���
^v���VO���j�n�7X\r�I�3�݊�sz#���]��P���gc�"���\���n��8�g���?���Eo����J���zv2�:�$��8P�Qyo%������D�Yr��h�-�i�Im�N_��SG��)���'�:���Rhhr�ذ(( �[����	��d��&�7�8���cߩ9�����QH�Q\=��K���d��$pza����s6>����/K���	.���[G �#�c�I�h�%����$��b�3y�+�+�G���Ԃ��$a�r���?^NkeY98ۨ�ŏ�]v�lNLK�d�A��?\�PM�6��ww���Ip'��ݝ�Np����5���K�{���W�Vm�L�>�Ǧ��`�T������(}����b���l�]�N����֜Ϋa&8t�/�I����+ᶾds�����3��[����
��;�;���N���+�̈�R�F��+�jx!�x�o< ĕ�H.Pp� -a��q�>��ۖ`�[�n-ը�,�_�w������;�9sa}�YN���hYٴo�̙9cN����y�/����R 
�ΝT�h����%�m�5T��Ei/��^��<��U�����b������&��~�7�g*X��L�P>��K�I��h��"��z}���_of;<��oC�X�Ar4�9���`jr2�|?��t�P�����|Ůx�mߊhÑ _NF�����\�����z����z'YA2ޥ�u��G1͹�T��R$P���M2u�V��	:}(oc,�R٣�]��a�x�T�B�q�n
9͈@�g�$�ݢu��]��=�����ݚ����T�'WU?���� �ې���.�6���>i�s���4bɚ�z�7��v�U�T" � 3�k(G�Ӿ��&�kn#���Y
��P����h;�w��G�t��� �E�탚)S����?G<���}���e�|�U❗t�	bҎkG�&�U
��<d���`�V<Jb@�%x�k�J�ɼ����A^���;)NH��7ӹl�k��ز.<}
����{� ���Vt�t�ק��󉇟
����_
w7ԾU5ѝvy���H��Ǘ����p腼��N���3� �
�h�X/��tw�4ެڿ��dG4�$k7?��~^t8!�[�L��a�k��"F�����B*0R�,��)Ȑ��Q�u�a��袲PY�R��t�@V 1S��'�(�vZr�L�N��-�o�g�,"�	�e�j��B�ۊ��Sۂ~0@͜�`8�M���>�Ha��E�eTßCg��K�[SA ���'�h�|Z�>8�omwۚL7i&�o��li��mn�z�>L&v(1�ʚ@:�R%�)c����l3��X��rũ���Gk�P���>>�YĦ_��T�@_�F.j9`����^�r@%�Q`��.��ѵ!���+M��\n�c���c&�ˠ^�R�/�$�C�� ��`\�ޣ�{���'��{}�ϐ������\{6�@-���8��|����>�*��������F�5���Ve�h(6ٹ�ĐY�&�@L���8���⨆~�\���.���aC��n�W�B��|26���l�ޞD�����%|>#������ rK�@cGs�x]iN�T6���FA��ɭ��O������E�������dn�ZsjMxV0���]�,Ґ�&����NU_&7a�ݢ��!�&����/�?^.�l�.8}\v���ˠ���ͥ� m��9,�5�Y;�CƦL��|T�#�(�����a��ڈ9<��{�4��eR;�~�);ZT3�ׯb���� �G
�u�3�Ɔ=�u� �r���]�k:�S�y�`�Z2Z�f~�_ێ�h�W���z��,O�Ý��Ew���̳������h�ڿ&�(�eO��gk-*Y!1��ٖ�R*҇F򰴔N
��_'�Y~����K]PR�_�#k�u*K��
yS�?_�f� �2H�x��{9�,"�6��gn����za��Br�)
���M���)�boD�uT�$�T4i�W1DBdt��~if62Ipj�MqB�x	�ټT�\&q�U��4�u�$��..�싮sH���?�AĜ_~I��{�q����V��Y��:r��v3�N�ufÿƒ_?��83Ctns6��=���}��S#�^��,#)fMb6T2��g�euI��Vev1�B�9�Ɵ����%`&ʎ\�Z��-.��,�M�~|���2M%T�1#����3d���g���dc����������Qq�ֹ��pi&!�:�M�r7��1A虌 Ƶ�Ý�����,l�j-���	�P����ǜ��:�Z��͓�<`�"w7�4�_;4n\T��q�yJi�	a(�n�3u�Xn?o��~�M�۝�\!\��jԿWm����}1�Yyk�ܭF�y�E�����Y��r��˟�b�&��(�84�����ZC�ǚ���bӟ�\�`����:���I���M��(_���V/��l2KTT�W�5�@$�(�h�OY���Q�*��J_�C�����MI$`�NDQ�NF�(si�߁Ȱ��,�/�Z���(*2����h��P��°�
��*ۇ�5���C^������@��A����:��q� �!�N��XK�ۅ��	��c�M9 �i!���M=F�mР�a��������Ba�@	��}��p�<��Ŷ���Q
�e�/��� 5ġIa[�cM�\N��
�t �������(?(��Q�/�+��O���0i�'&n�`�bV�]� 6oG�g�oH���l� g���3BE�jq#ږ�����u1�+�1'�p�`���7/��dP:��t�tX?�Qw8�W>�7���K cW���2	�� �Yy�)�q<z�.^�aL�$�G��ԙ�W0R���!@��W�<64���4���(^�Tg�x8�W#���S� d���W"я :M�� �2͹�%��ۄ<tX�x�v�z6�5�� n��$��7�Ǻh57�`h�����v�j�A����q�q3��nY,� ��rc7�jU=A��-:�36y��9�j�Yxy�"q7��0��0��98�����DN���\n�׋��y^T��⁐��)�@�٣�h�����������'�Z�Mqi����P~�N���n��}�9�����@�b�|���rQ��/�fs�qa�ys��L�3F��P�b�[�%{��N�}����z�XY��;��E���{��q���&(��O��MV`FD�޶�{o�2l��xN����x�O�6<�uU��{�����e˟��Ou>'p��}�`9Jiy>=���Z����"!߸����#��D�⿝����m����h1>%�a�ޟ��6�$C;�ھ�� 7P
'8v0m</J�^�W�#'��K�å�X:��o-��Am�5 q1f@�����V���A���Ⅽf� W��'���53V�pX�j[�ǚ�y�H;��(� �!Iwk��4
��ԙ�`bB��}a�����6���]���κ��KM硜�%T��d��u
*k��`ط����Bt�Cy^GlYY�;ᯏ�/oG.O�g�G��N�2��@�'���CG��zn��u͏.ô�]R)�˦�����eca]Q�]�X?��Q��;oJ�.6� Tcr��V�/��t��YU	�Xe��jq��O�ᯞ��yY�0ga����������
�h7QA�Y�-%���!��.7�#�[�\���8�8^P��c۠T�8Ý��d*�T�����ݖ!��\��b�H��}�1^^��U?݆�ubr��`Z_����c��-�m�O�!
�Еￕ*cA�f��QKs'f�[y-�R��> ��Ç	2�U�5�c��~���b��|�)�G�L�����h���-X!�ƒ2n�0{��?$�s���z?'��i�XX]狂��6��e�]�:�.^7�f?lB�p6Z��6(��O�y�)�Ο��f�����p�Ѿ���{��A��Vd�VIvB�%/9i��;鮽t�p�GQ�L���/�)SR5[�������]��Q��S`���S&��뀫����b�5�%�"bMض�Q܁���E���ع��Q���id�!mr�ag}D���X���k��x���?�d�}%�>��"T7�r�A���N���χ�SUG�X~�q�T;�y8xrySD0u��ZG��6}]�=��P�ӳ�+�����;�Dux+	���l_��!
�3������.?W5=+�\�t�6q[��N�9���?�0���v���v?���j��h���j���j�߈�`�W�.stf�/y|�Aq*R�/�'G���9<v��Y��Fi�6�;��&"5;=Н=���_��wژ�	nV�`�'#�O'�VY��߮ZUA�ŌQy|�hu���Z�h�o2����j�N��4�� @��o���&e���'�����}x��b��ꞓ�LPw*^����L�):i���M����;]*�u�$��*3z�7.M�O�ȹS U8Y )2����)O��x�f�E�2+���k��ꔄ^]��ݡE���K�U�&��=� ~J���u���5c���^���ӂJ���6�	����I/<�;+]G�6�Wmq�ko �_s��/��E9���<6NZR'��@ax��ǟEK5Ê�y���dO.������~X�IZď�n��Q����r��;�v�M�{8��͜Ų��1/�K�p����$�痀UY�S��_XL�Ȓ49�zY0����6���F�P$����2��ƛ�QN��Y$/���^l'L�l����^Z�N���	�~
��|#���r!<[ja}|�NV.�ˊ�H��SD���MT�:e�0�O��4&W���]j�^zf>���c�˘������6�( �i�mp#3(��&�O����̈��l)�P����DK�b���
鱃��=��ND�tc>T$��j&{�f4��jB׶�!Kp�����>�Z��v�4sʛ�Zz~ځ:�Y�Q�}��`�|��%�0�9�5���ȷ�d�{Tp�괕j����d�P�.^5]z0#6a�;(xBw�#ͷ&\u"��ڡe�Y��Hg������44�	Z���*I�/�x��%N��傢�w�'����i��	�;�AT^s~�����h�F�Kp��ٸv������GX�%;i�
�ڵ��\ �����]�VP����+��e���l��ͺ�ł�b� �g�
�	m*h����e��sTG&r��-�F�Bĺ%�|5��w��P[�HEJ����ƻzwHU����K�x;�g!�Ì*��ݑ��N���|��h�׬�jB�ྃ���i��3�{q'���o6}��r�,��Q��[jj��*��M�%ԁ�E����� ���C�Ksر5��9Fӻ��He��ޓ��hu�k��bo�͛���|�щ7�.JK�d��N����8����f�H�.�f�B�[/����,Ka(�Bz¯�m5���8ۿY�n�"��&�j]3�k&�b���J�J�W�<Y�%eyI'�3o�$��e�L\�iD1$�}�y����tC>e����k�%:��؇ƴ���_�����ݘ��X>Ƴ��&����r����(��]�^��p����X*�y�.�Ω�q��W�����xE�����W�T"��?��BxT/����d^�x�b�% A	�����`�LA���ب��d��N�DE�\����`��0S�Qf�ƍ�cX��(|���G����U+s��u˾�\F���y7���3WE�]���0�d�gu�M.��J���F�}�J�>��(Y��?=�<��W�����j�ޅ��#�0l~�떜^uPTn��V�
�^��y����]D��o/1���;��Y|���/���I��(q��^��ZGp!/h=��ͬj+�~Z�B�TO�|y�c)Ops��p�%�:�M����%��;��ͫ�L�֔5d�L�������|,|�꩷Fc�!H��/\ډ�7C�̈ǜ��Y���ﱅr��'�ԯ��q�ycl-��?�~2��<���3P��;�whUµYĴ�]E����B�١mM�g+���Wu"�u)l��=Lee�yX9z��##sEY�Lӟ�-���~��54z�c0� z������Ji�����fi������jn��?��$PPz�6t�ĻUO��/����^����׮bMz���ܭ�N���U�fF���i,�.�$�Z��
<�F?�����o��-���}O��퀘嵭�����k�]���6��w��؉��+|^�QCe'M�S�>e2#vі;o��}'c�n�]5�����;1C���^����`�l	T����4mm�؆.mK{
��������I���� �}GHy��r���|9A���N�[
ݳ��8����K��2�e�ڄ�<P�.*�xb�W����Vr���S����]�|k>�r)��Ţ�r�x��.<?̍?��'�x�jƌ��e ����~��I��"�o�H�8.'���۶�����u���c�t�pү�ɐ*��S���;��l�}���lF�+���l�]A��۔�\����۩�_��QVD�������t�Xלs<�/��<�,����Y�~��>xT�����Q��_Oxm/M�����Z����&$����FF�0+�[Nz�7	T�Xv��(X��O�,�3��,=/i����T��xM򺡵XߙTd~-Y~��	��}����uR�
��p�����kl�9�U6�̌x^���-��{>X�Z��Wq4ѸЧ��u�jс���;�E������x��Mh��__
Kz'�,c��wrZ"�`�6�Ƴ7peZ�o�tdeȄ/hkJa�KT~�6�o���7�������ڻ����`�ɿ���J�9������ۅ��۔e1����9-���1���y}�1y-�5����e��e��4���I�C�@��yo�"��G�"��i��O����ҥ\4�ٿָpXN`>�@B/hH3D�.���}r;�5��	��aK��X�Y+ ��*���i1�ݗz�qĮz�8���Tp���n�,��'*�O(T�K\u�
D��%�H4�njuu�֔mU�,r�g۟��Y,��hO�;�B6M_^b�t�g!��;�P��-�z���$�.,>������x*�jzpsD2��T�C���Y:�y��@kUȒ���:��k˹���zd)��ok��t�yW
,.�v���|���ꌐ�����+m[À��*��I����"	�������ލ9�/.;�9R��JӔ�Y㣨�a`+MuyS?|2B�i�9|�K_���XLZe��F����~e�2X)�1mª�b��;����Vg�	]�S8	r�/St��,H��T�e"��-�56W�
��7/��o��[�$�U�(F}\�bL�B���
<B��K!��g���,���-i\� ��!�Jcq�T �w�Ŀ�?�!��\���CCi�Z�,�r�)S�<�����in��P�zw��|�}͈),O6����,�~y0��H������^*���� g
gƑO{2P-����<nЌ�ա������5 Uk���3;GFY$�����7�%!M�h�5�ܗ�5��{LT�*&��Lw�7�&pj�}�ͳ��?�x8�)����-�L����ū���8�j��a�=C�xT+���~� i83J1����)�ҳK� @|��M��I@	�fA��r����S5gHN��z����D��)���0�z
��Q�q*(�D?���~�lV�O��7O�=��K�v[�$����L~�Y�1@D35@}��'��7���? )j����fp��kh��a�Bu��`�<��Iv�����
^>����Kވ򌦗R��1Y�G�T����H�[��Q��~ڵ�d�"�Mh�S�>��cŦ�eE��S7�D��F��+��,�������bie*��?�-�;vw|3�@vO������_�=윲��@��,.=�q�oh���9%I��W�p��w�`�2?��,���^u��.�Bʕ?���n]S�����(�7�G%I��c(�[�Q1�Z��u{{�G�Ν�`[m)(��A̿�&'0��D�����A�+g3O (L����t�V{=����S�d�-,L�h�f���V^�0��V$8�=g�Bt�M�e����?���޳R������>�J�mF����q�Z��n��Q�P6
�<+�{d@ÑF������%�H[�PeW9�'#���]�%�3��c~��&-�S��6�s�A�}9;'�����kr���U����
�0��n71R&��U�TN8����A�ԁ��Y�e<�'��`*�SF��FC.�:e��<��<nd����D����yB��1U�d:�J	�BZ[]>M G��`�z��r�����K�������ҦoW�Ar�m�烱>7p�[��X}����R1��0D~kU
c�C��Y+�����l_M$�Yw4:֙�5��)�Z���A��21c(�`�V�I�5�K^�%�6|��P(S�q�}�-�h6UУ%/G��b6�o���B�z�WA�����&����x�|]�\:��C��Y���ڣ�v�R�B�}k �����:B9Q�C#�v�LnP97K
���ڐ'���	��H� �XL�i�ao��!��}z�,�GK�=��:��3�� �['T��I��
����i�ې���1���PDq'w�@t��1���	����O����Q_�
��%<8��1q͌a�g[�#ƀ�X��ԧ����tE.XCW2��/w2���d_�"E���|�EeNg� �D�ŽD\���]t�!�������]J��Э�j9��u�CK�]��|����
6J��}�m�$-��m�yM%uBT(��6Mtn{܃�XZw�7?���i��)�֎/wBx�p޺�0H-4I��b2�kOI��/�N*\��?���Ew�NB $�`�-Q-�����f��c'j��O�r�+�U�3sj��zT#�5٪�P��Ũ�Å��S��v���*_܎����AN�P3�����l�%ku�]=_;��$�
���z �A�Cn45�� �ǃ�|#*�����J@Ir�O�"��Z�Ѳ���dKC�I某�%�p/|�žJc�L|?u!�� 7�j�	B{Wx>S&g�ɟ��1��#{w�2�c2�-���(�Yy�_X��s����t�jL����0$(�0���5?^4x�M��J��j�})}=cH���kCdK$�-w"�	r�ñv�]j[Bb/�z��Vg̲���8�L�ispk�¦n�L�8)�����h���J ʅ�4��")H�eHX��l��m����L�e������Ӻ�s0��������7�\�B7��
F�C*hރ�����PCg�����]3(����ǉ��8��r2�ڕ�B��bV���6DT�/�=�+�V&NV��@���w��.� �C�Nn��Pִ�b���=L�sZv&����@����C���݉E��d�g?*����"z�K��xg�Î�%��T݅��Ϣ�~ ܎1�/��s�4��ٺ#n��\�G��W.���߱�"��e&'@�Y�Gf'F+�����0������(�gr9�T�Gm�;�{�fG.c�\�N�"j�nn�%!f�������2T3�!0�8��=���Ϛ#tbq58О9c,"5QqbA�S_4'D�M�{!���>�#�8Z�rWn6�<3�]��{��Gf�;|�b���'Fڷ��CB�%���Ɇ�5ﵵ�y��υ�De!n�J#�~��%P�D5��o�� ����g�,f��Qq�Z�t�_��d*���EX8��KhN���K=
\Ծ/s#��#ip^?�������B�G ��(���:xܕ`�:`:v�.��A.��_+S\�a)<�Q��Ԅ��\CG/�}�ق��9�Wf�)"L��� ܲ�X��/��*%TޝZq�߱
@�dq�?ŗm���#��@<�Z��k�kw�g�I(��4>[mݱ����%anY�r}V�V٧���K��@���U�����C��]
D3E��7��T���V���2GBԎ��[86�A�V���..�n�������x�S {-�DG,2��VM�| Mu&����*ȑ��H}�u�n���=&ꐂD�@��ba�K�M"�?a�S���P����0�v�)�w�l)	��a��)�0���u�����K����9�ޮ?|:��U}�x8��}N)���_����D��$��c�|�vzp/��j>��o�[*7R�*�5rT0ᴝ�.�?믔���3V�*����%8VUJ����f���9"�oz�s3m�j���� �{�����������	nI,G���98��fG ,��;�AgMP�=��U��<R'���!�Aȫ�SZv̩�ԔI���1`�l�~h-@s|��R�N�j �C
S�tW ��h�oD��D�=�m�����xz�gơF�"}�G�z��A�|6���R��ۺ�O �wEۘ��_�����i�n PL�&���R�^�=��?�*j~@"	0�UV�WB�6ħ}+����)�b_8�6�� \r���>��v����,y��%'n�W��z(kh@(��ť]�{�'��g��I��j<A		}����`�u�S��Mn3����s��&�E05MӰS#�F#�YLxdi�i�s�#�w�|z�0�&7�NPA�5Žߤ�����qy��k��}������2UtV�J���֣V�d�U6������˔������.���2�Ƕ#7�c��EO!ӛnlkty��k@`]�q�d2fF��(}����ʡWxu��O���EjyӃ�|
���R�P�%o'�Eܝ���}��{v��1a���}��P���(�W�Կ�۪�Ѝ�ܖsmM�q����$��V}�Z����c���Ыv��P���\(q�L�W��U;/Kq}�����vb��#���3ި�Y$A����+�U�򜣆�����P��7j+���Z`*?G]�;�V�!%�{p�ޭc�]AA1*�ڍ�op�՛��+����!7xD�<�w1޵�p��K��z�����.0
=�7&{H��n��IS��s���=/g۽r��8���������.vC�и#�	���+[�=��jqC��(�#3:�aB�B�����Vj&����6��^&QM�T�ϥ"b����Yg1T5T�Ŕ8XO�EP��m��b��r�)O	6��X!����A\Y�6�f�(��k�Y�a�oY��"�M�X~�Z!���}�w�	n�V'��� �r\��Z7����vzƴ)!��6��aN�L�N��zI~�����z��ٯ�ub���fDaBX��;C�@���-�f�^sbw�ۇS[,�ޚ!-%��5O$����,j�y��#Pn����#��0�K�$�Go]n�]gi�}o �*4�ܟ�I���S���c�88�]�4���L��	��?�|)B�q��*5Ǝ���b �JUR`���]]�7��[_Β��!�)��4��������w�s���*8���m�b9����������K��W��kl�ڞ��=�ia�X����tfkjB������u�����y2L��cߣ�uZ��'i�e҃�r���f�~K��a}��5(��H�����w�3���!�H#2?L�&T��rw�p�Q��LBB8PKݤ�L#��
�Bf}�Y���˷��A|1�4�mw��w�:ѷD�g��͑�.7�������Kn/Ab���a��)5J\P%8e��c�d닯@�.�2 �]���8g4n=N(J��\�]s$\|I�<��B����\J���"G0�ln։v18���s&�^��������ڄ� Ot9w"9n��苽���c�Oޚ���Cu� c�v�B8&B�0!ב9��~��^��_�q�Z9�ü�6HY�2Z�Z8��:,'м�q4�d������)z�"���W^��C��(������o_[��E3�uiב�k���A>B���v�R����i��Җ�װ}�6~���u�����:�OG8cwtQ��\�T={ʬ���>���D?����3Ӳ�:A/+�q���֭j�\���a�t�n�z
�L��Fi��O����kԃ����������AL�E������nO�ܑ=��ҕ���u݆`����,��yǝh�G���:P$H�T�,��hr	��>P1�j���тe(���F�x)��x-�N�{��~R� @K$�sR0�MJ�8�ǆ�@7e��c�"��LØ� �.�k����@��Y9�&%@����w����:��S������]Xkt�Xl��:"�<�<�z���}�vdd:��nl�Om��2�v�E����<����eGh�u)Ռ�����n����R�w-�w�%��RJ�䲥\�|���x�W_u���o�;W�4��� ˃� (���	��ghG��@�]P�����z�2�8=��xyW�?�R<95�[�+ڋ����_��s���q�}z4q� X	��5TP���������	�q���F��1����K�+	A�q������͛�0S��1C@���5^9�T#��ۇ$���!���3���s���8tn:�v�k����˴r"��ͧ���ϊy%;��,���ozB��D1n:K�L���N����b�q����-Y�EP�#��1w�=O��Of�u+)���n����ǎ8�=����_S��r����,�Ӳ.��:Oڝ�m���F�I,c�@�|�$4%I�����`U1���׻t��|�ھ+�̥=�@&<2��v�/:���| ����^�3����; ]ͪ��<�b����3���^�����xL�`d�r��c:�9Wg9ƥ��FQ��M�	NB��~+�����ig�;�-Sj&��^�x�}n2(���=;�(�v�%^o��X�$����S��=��7��@.ݜ��RL���m�jG+z ��i�Х�$\�B7����s�@���5�׌��|3��G����,���>R�^����ł�A�*gh;�S�iP>�KCy\3��q�Y �2��T�@��}�a_�!ۛ�t/��<�ܝ�:滄s
iLn5��-5��FP�v#�HN�I� �����Vxw��i�`��²<�'�+��m�EÚB�<9b�ऑ�c����`yW��"/���$�β�Z<v��.�mVX��A%!REk�n@2�Ab"A�#�<��2^�^[��d ���O������ڸQĶ�UΛ��	���p�ݼv��������0����B+���F9Ll�8L�6����#32��oU_A�
�w�1�m�04$��;�篞v�GP �'V|3rp�����^�*��16�_�!����5�%�t���+~",���pQ�g3�ytE�E�"'�\�Ѹ#�A��qю6dJ��K؜Y�-LTgꧣ��)j�Q�/㱣f��}�
�_�o�z��ۘG
�u�dĹ�β���bێ��wo�Ce+�O#�������>�͍�Y+Z@�nB��$yL�-�FM��|��D>@�F�O���bW�ڔ�g��)�.[�ZF�.��7nù
��|%�p��9�vz�>���V7ӵ$��t�������ɀ���ψ���2y7MY�!�((����'�曅 �����t�����y���eE� 9����*>�R�M.�-�B#Kа��i��d�y*�Đj�b$���
���|3aF��G�l8��@�{j��z&X*� ��[9��P��
��~/�/��<�� HL���W�9X����<P�P�������.q��G@�I�jr\���|���n��j��?��1�V'}�C
�C@�1=��06��
����W�v*e�;҂з��-pr�i�;�o5��ey}���-�>@T�k�p����
����V?�ّ����124A��ڣ7y�ە	��c` T	3&��!��G�#��p<���P�������M}Iq $���f�*�6C$-����O��`�OܜI�vyk��tc��+��ܸ�X�v�����+�ҒR}A���1,�8'����T��?(�~Z_K�j�����X	p;
k �>�ǕږlL��0�j;���Q[8����G�2������ S��NAVR�<�����
����y�7n�5c��+W4<��b�ٌ�=mK� ��0�ҴЂ��BR���_�T��>б�a�X��Qg�괔���Db�K�@<3l���6T����YQ�2	��g��ĥ��K
���v:�g:~����j�l5�>C5�ﳬ�����oij��Rl�l�i�p�y��L����^���}�L���d�Ӏ<7~��b�<Y���t�xT
��uC-�Y:y�QT�<�X�`��7/�L��d�?�GXL�|f	p���P��m���z�7�VfҸ�b�=���c���`_��xr��H�po�+l���i���ޚ���XH=�C�_t��D�cP����.�BMM�J�����aO���,3�+
��7YW�F0L4gn��;��
c
n-0*��xTC3	f���I�x �=m��\�|�� l&J���/v������֗������>�a��/���2��A���jВ��
~ �F�8��h~�C>8mu�a���t�Y~Q�q8nPq��A���	�G���A�hŊ91��;�����~(���:F[���^ۯ�A(*~��CЁ`3��3-����u�Et��kA���I:�C�wE@��m�vaiv��:gv<	�vFu���8k;�ݹF�u��c���GV�iJ��v��a�e��?��aM���0��ޛ���iV����
�zh�U���SUQ�5���b8�P���Ga�l��@菕��=�a�T]=��r���3awww��f�g���;�Ƣ����:������b�>3����g,n�hʆ<nԇ;ԉ�;����q���/	2�̰P9^���5�Y��A<� ���wA�,���6����/�74>O39�5��0$^|ߨ�y)>o���E���f�'��ۨ�bZ�h��C���{r��P�� ���b�yl��{�^�� >��7�ׅ�����f��qes�G%p��mGp �6v�TYY��M�������dw��|J�!')��|�zP[�����d��/)y�诣���DE�_F��R6~:����`���CU�m�Ŀx��.O�'��B���>J�]�]<�ĖO��J�	��f�kJ�E;�i�� 	�W��B/��D_�x�.Z�km7��۵��rVI���\U`�(�O���|�[��/6EV=�+��v��%���ܢ8`L�+�#BR�1zZ �"T�I~q��8!�5V��pi��38q��T�Z��Dr)���Q���s���܃�+m^\yt-×�lT�ч�3�|ot8ZR5�bn	2�%`��04�d�aB^4��{���U�T�Y�,�E�S�P?�/G�&��iq���j��	C$H�!*��s?P2Wr2vr�n3��C��SX���A�ik��F0�R�� ���)����G�Oh͑b�&��k��ς��E���Hg��H8
O��Y��a@��� ��j���C` �B��TJ�%��I���$�q�Oh�K
���?!��Nh�?�B�����{��܅d��Z��-
+#q �y�s�Phm���a)�`?��y�?��OB�lSޏ���s�&*}�5t�w��"��?�AS$�!���|�i������[D�jw����?6���UW�̟���k�L�`�����CR�[42h�h���Cⶅ?�R��2�5$��!3����ꚊH��G��(&�&��j�'f�)#K�-�&!���B��p�8P�~l�����~� u�"r��\�ȝ���z�B��7��JU	���5'�v�[ag��ߠ����
Q� �A�4�R�!'i�Qg�p�� Ɏԇz�N`i��Y�d�Kի�Iq'�P���M��Wq5�EC�P ����H�
�C/Ifx9�ǒ,V?@���=�?J-�\�>ް"�b�'� ���5�(���c=)zڪߢs�A�̜t�(XQ�4H�Ұ�����2��-� �=DtRf60K������#�}H
�M]i�/��|���߫�������n]iW�}�	_��t���,l��b�= c�+/L��0�!,K�� �� �H*��hPj����J_���s����M:�&ް�[0��A�x ů��6V�ǩ�7���Ö;�o/ w��/2��#�#��)����%W:��$5I1��(j�!���Q�@��$�u=��?���j����u����\l �o���l�+�
������T1�� ���ΰ���Z��[���_]�v���o�3��z���(*�@�L]%a7vR��*�;���7K;��}�ӹ��~)�R�c��[�W�WB�4[f�'��*QE�q�[�(wȮ���#�ז=�������v�7��TV�����:@�����(df��ޔ��Y{���๸~��p�z�y��+�avG�4�U���!��-����j�]��dg�>�B�Sbu�=>ڠ�>\��j1PY}���2u��;#u�쑞��<�:�x���q�:���l�Wj%R�{x[�^�ȃ�A�n�Dl�|��<��%O��\��u���6I���8$!��L�J�щ����u�_����o�}#<}}& )G�òT�H�q����ڞ��|2R�]�3�!��|����g����(Dc���!�	��q�ߗ�h���N�t�/�'�����EB�� �I�����&�T�5�(f���P��"�B4Ht��P�:25��ȅj�#�M�~�^��ܱ(��NC*��N-S5�&����;�m�������f��[w.�~~p�(�����ŏ�����3��A�;l�x�{Ux�zg�\ʱ�%�g ���}�O6��B���M_�?Q�������[t0
����PT4a�hڔ���������oF�2rrv�ԛ�㯅^�q���Ǔ�����j��ڼ	��t�HE�ނҫ�J��(@jD�H(]@�H��.U�-�*z��]��7�f��53��䞳���쳟��uW��E<��J%�И����rC%6dA��{�f��1�E�5m���_ד��Y�7�����)��B]g�O�b/��)���yy�&�4bƋ~U�Hs��uE��inl(���L�jt��`��N��ht��n�P����W���a�雥w�~�JV:���m;%�mB"���R ��{=߾�,���r����7����c�V�,kC�rw(*�e���#���v�F֜�
���^	��g�?:bu��;&Ism�U�f�Tf�fZ|�]ay X�3����>���޹���Ns<�H�d�@�m�s��Ϻ>���|�~���i�5%�s�hc�k?T�v���eH�N\�0ְ�[�im������6L�!�$,Z��ɋ�f�V06}��S	��3�,�q',���:��jģ��#���J��?j>3��_B��t��*�h1{�yI	���T�ߏ��2�kJ�"�\O������_�81r�k>=X}�C�)��>J\g�	H-2L��#�`�V�IǟCIqd����!��6����x�X1�8�*���1�dE� ���^���X�J�"��p-�N^��*��%l�_��ʇeo�^�to2<�����uRVs����\�[qO���m�̗��>>2ҿ���P�g>�&�(�_���d�/�Y��0ik	g���)�
<<c���A᎟-��L�����_{��tv�����;�/R%{��^��ף>�U��W�,���"�3d�{�²�?,9�5�Ɏ��
�O��̴�&j�[/�J~���ݏd�-2"�ʌL��#���X\��~�M�W�-r�#࣏Qq���VT"զ���d���h�R9@R���ё��ExDu�u�?�ѠN��9f-''��>�6��Bt z��ӫ�(�
��틮Y�AKE���.���鞲֡��@k�U?V�Zd1�2�$wW�-d�@&�A�\���A���hSI'T��C�x����&�NN������IE4V��J��JD�Pxj�7�8�^[�t���%:��!Q;NO����;��@��X�FQ {�-�w]p8ִ"�f��[mS�jW�l��Y��#��4O�����j��
��g^T�s�Ʋr�u0��7�\�Օs?|��u��������f5�Qt�E���OP^O+TY�k{~4�|
�#㝬��M����p~��HT�e�_��V4����'��g\N���J�|��do���*pNnnL'038GR㆖�s��o������������+/(Rh��z��Z67_21���6��5X�̙�݁�#�y�@D���P1���@���� ���%��a�D	Gwd�EX�)�1�/SMw;�>��Ԋ���=LS��[��P+ d�95� ����Ŭ��z�k�U9'�0KY�hW �Z).Z_��?�h-�D
�BRr��L���q���n:G˦*"���
XSu���%�����nB����o������_�#Da>�A����(h��e��J\,��E��"�ח�>0+��o �#�[�q��B9�Z������ 0䥮W�*�!����;Z��@�:�O�@P�m��y�0� l�#�/�0U�DH�Y�E�_t.#?T{Z�V�L֗��9�1*��;i�0�m�����'�̽�<v�T�ޢ���/4Є�Z���J��Vkf9����FI�T�ԙ]Q�0B��N���{!�6q�vƻ�
��O��C�R8�����Z�	�Hۗ�u|����"BZ頚r��i�v����ɩ�&���`��:c���mK�0 �},��ϖ�8m�|����a�ʳ�'q��$�W�RG2��&���;�|}��� ����r6��J �X�2$�����R<���!V�a��PI���{M�Fu�٫�04��+�\��7� �_Ri����*u����'�Y�,���"�Yp��p~��6vvvi))���S6�2>Lm�w�2���)����2�2R����<S'H�T�d�
lsC5�4��?<�6���`?+�4�(X_�[�l�k�iZq�Jz�V;!z&�+�����m-�2Rl=a����𺵦'S��9R��btuQ�t��9�/u|"lgR'�Z���_�±�+V�8�D�h%\W��乚&�7�mJ$���;#y��O�z^x_ 8��y{���ADa������.��x=���D_��*+T���07�5e:��>N��(�][�˾8��ୗ;D��0�����Y�8����[�˞9�����q��G���b�ǡ��2t6�<т��`����x���v�>R)�k����'���/����#d={��m�Y	~�b#t�h,��.NK�V�+y�YC��.w�NYT�kI��>��E�)�-�gJ�.Q��B:BHG7��n�s�����/^�s�].��;�@�Ҳ��g����Lwr�H}	�1�� 9fC
}@5�}��i^C�^�V���q�#�9�U��a��~�O?�
jw���\��&%��z�	�`�$' u��:�k.^�׹��{��>�_wڦ#*���_��g-Q~Q�2��E������z�m������"�$�S�|�E?�h\���1�z*���.�c]?\]s:k�J�/,P���S3�_�����_�ƪrEB��K��}&sR� )i�Fx-q��N=D����!AEت�il5�Fh�=�[͜/`�k®�xX
���7�0c>-�{��L���[��m;s�S���RHŠYg{�۷��0�������t?�6�n ���X5U����&���n<��u�r�JH3ou�˭wM��r��%<=+7�C�ۮ�Q����rj��T�|��Y)�N���*z���Wz��Ol�}�~6��W�L�2�{����j���(�d�HY0N� ����C�ng"�Ķ��iХ����j*��ZFfl�	�C_��n��A�6�"$5��!�K�1�z��)�;z%�^qj����b�w=��d�W9]��<N��.�,Y�?N�n.������O�"��3�fl�B����.�2*$���T�g̕/�v_J��?�jI,[e��{w-kǿ�p`���t��H�ÖN�p�m�g9܂-F��2��8�b�M��� �ꛗb���չW�'5ԛ�NW�P�̖y��&j����p�7��p85���[r��$8�֔~0NC���H��k쫇a|�yee�1����'F�]+"�x#��zJir��b�u�CS@06��4u�*Y+�	.��'��ƦE�VO����^]�*C�{2#cS<X�Ɔ�j����w&s���Vz��eE�R6X��F5�g�BU�t)۔}��0{�)�&p�,WEP�tɧ���MV$�΍�2u�8�������\��;�1��𫡌f�J� =�ɒ��w3���W;�M�b�*)��H��W~�V�I�5�O�{���;qx��o��P��锃"����	�A���Ch��*�w�Zݭ�^�O\��dx�i5�;ٛo�ہ�q_����Ę�N{�;���h�W.V0�x��"�v*��ʹO�5n�������Y��	/Y,��7���ke��A��ƎW�]�7��/��)f�Z�X	��ɭ��5�"�j����Ki��fY2D5�ۯTm<v��&=ӝA�m����cU���y#�c��8�O{�^w $��l{�@Hh��0�o�k>و~����2gH+[YY=m!��}n��m�7��F[6�D
�Gp�k�/�Z����ܳ��YJr���8U����rwj�b=cyw�i�����qc�˾��?Dpu2��JC��M.��ޭcA惱�ic0_����+�_���b\g6��:_SC.�,���!Q�]''��i�#��n����>i%���L�%-A4�����V^'L��<"\��saw탹��_��>/,^Y`�:��069���Zu�5;[AA��<X�#:��<s�������#c�����W^R���~uV%�O!
�j��K]$�>i�d�U?z^�����Y=�[N�RP�?ٞ���޾�>:�w�Jq�i��	�\b�����������[bbLKU`1`�v��[��z�ּ��\���N3�f�������sۛ����k��V�_(���N�a/i�~mZ��^h�x ���;�7�[��(�4���s�����M�;�g>n���舎�6��(�0���Q,>�/l�HP��!��3ȁ��� 1��}�Oӕ������L�Sp�w��چΩ��HK��r~�_��{tyZ�`�5f���Kw,�(��<C-�ߺ��.:�Ye̲C����D��$Q]^Y1��(�r���Jng��m�"�5�������ۘ�W0�Ǆ��{���_cA��G��xm��g��M{�n��o�6m��ķǊ�o�$�:e~�.6m�k�8f��g�����T��"�U�&�I7,��t��M�n��C�񍤢߷��'���ȘE(���}���jK3L�rk���A��D@���ag�<eD::J�9.]z���%W�֒�O�H�̘�1餛a;�^����5*�W�I'����JR#9�@W86��tz1�B��!��H�9:.�R�`�+���n���L��r8>"G�!��Ǐ2����F�`]�]gQ�4����ɻk�$��o۟X����{�L���./��~���ߙl
�%�������?8`D
l�I։���Yg�8�����RF��U�8�ň���{M�z�6y�vZ��b�X��;e:)I���?=��o���eⳁ��3(�Ţ�$��{��K,W��fw�d���v��@���g�B�s�㙂�tl<QT@;�~7gw�������V����;�� ���lHK���,�TΘ��f, m������,�=f��y����	�I�m����ӂ��Cb��	\?��E����_��ֿ��.{��������Pq/5.�����Z-G?EQ�	1�%�@ �0�):~�w��d�h��#f��Y��4���<fox�D������b�V�"E������&o�E���jT�b\Z������r�]32���E��-�BCp�������&�E<Id}���"Ƴ���6lT��K�z�ļ���;�4�7n\|��[�J�lp���!�AD�x��0Τ/K��歭�­:�8�+]���ɼ���J�Q 2��]��~��
�)���x�`��D�00��8���/p��^��q�ڲNu��[��{-�2��E�j��y��U�J$<+ #�VW=�q�&�Z��Y �6[�{U.Hd����%kve1���.�,z^������%�'���O��7c���H�+��·}��㶞
��ށ˖hj�ӄ#��.o֯tZR|�k�/��)#y�f��'�H@fXs��n�Ш"V��m��*�U�ٌ�~�p',����~:�\?��P���������\+p�gkP���
@�Z	��;��Ջ���@(����d::���)�R/�v��F�6m'\ھGt�q\���3�;��~�0�Dt�ot��t�ԁ���ͯ��q�r�p�M�H�g��d�~���Jf�/#/���a��ebhg;.�N��r��͠���p��޻�$.ζ��NR0\;�hbi�>��T['B���Є"�6!M�SS`��~�(����z(̋�)�Q����D,7G����`���o��JUN�GƦ��`;S�/XOqY|=gr-ѻ�N��!!*qz5�^k��9ĩ[#3(Ʉ[�8�����?b��K�<Q�$Ԟ:B�n��2�Mv�y����c%R�nL�y
�5Z��w�/菑��!/�7*y0���*�:�]������rtŚh$��ܸ�I`N
�K�n֍�t{ᒧ�e2�����K6NrzM;@�-*��ǭb`y�^�G_��[�_�7jj��1B��c���N0�V	���b/A%^9���y	�r�}`�t�w!�C&�|L�y����ߕ*Я:j�O�@0rF������(��R$�dg���x��S�A>���ڄ��y��������:Ij�ih���c���:hJ��Dm��G\���3�=�F��?b�����������Q��d7:XxCj���9N������(�H�-�%���?x�S��^���< eK��q3�%�e�(+��P>=zs�E�7Y������,�P��P�Y�*��2J�~��DaT�=Yb�m�ű��������� �(6Q«�י?�싴yް�[�˒Q��<ojoh���P���o,����!x��E��k�o1s�n���m�&ry��;s�KZ��"P׶���2UK�7,��.�~�&˫�I qs�QOV�����)�F������;���51���[�G�������6��Џ?��i�W�~/��%������~�,�6pus���fY�	:"�jl�7���7ǈͻ��G�������.���ً���<����`ff@�����!�G[!��� �t�lοi�إ��C�8e�6��g+G "�� N��W��d ��i 0 `M���i�E����n�mԄ .g���w�e�� � ��u����3 �\�Nˑ!�/{ĭ3S@3/�T�T�~������`�E0fi�ׁ�~�гF�6ZV ����|h��xuۙ��; x?S�n�O+d�%hX(�U �
=��]�A���b�
���W���+��
`y��%7�؉������"H��\���V_pOCf���JNoK�!��ED�Q��2�j��z��w�h�|��O�ue�և·�=?[�UC�R�r�=�a��+�.'

�Oߧ�A�>�������+&�����D�C�+1�\֩%�������ww�G���G>���_og���������;��D�큸����������޳����U�n?�/PK   �C]YC��cx  ��  /   images/92d0aaf4-7c05-4843-a3a7-a4d3b320fab8.png�TS��/�4� M�"��B�Tz�H �PD� D����B��%����"(�y�����rg�{�̬5g-4��g?���r�{�M�,�,z�P�*B��@謘��tT;�������s�G�8�	���ͭqֈK��>Xig7�t0�rp�k�:�z!q�.H����Jc�� �MC�J!���A�І!~H�s�/W7a�������s�b��U�5���
><����!�u� h��,���T���r���TR�vQr��\]�U$�e�a2�J2rp)9yUUY��_�0���zUW�/q�NC������I)H��y�ȩ��������K
)��8�`)o��s�E����}qho��{g� �����V`}�a�������d��}e�ee�&ts���7��p7W$�Ez����?��(��?��?`����  h�@��`��P���q�9���_��U��O��+R/�y�߶_E��_���ٌC��{V��������`�R_U?�3������7|.��&A+����H˩H�J�
ʻ��+]����9RP��E��?�.��>�)%�"%3�WPU��*�[���쟤7����TQ|�WR�s7g��I�����u!Bc�=�2���^U���.
�F T/z�㜽]�u5��i4�M���U�M�)����&SQ�K�(�)I��U\�ar���.����q8����?O���+��oR�ݐ�*npY)y������U�Y�YA
�"�tSts�C*�������3�_�h�8��9�*���I�]a�R0�2�J��R������e�J��0��������_�P�	�롊�,�d������"��uo4p��������Ho��pEEſ�_F#1ֺh`��L��r��d�/Kʊ���O7��,o��L̐����A�qU�]������	������m�B!��S��I���r�Cjy /�w��d��s�n��\Q�M���&S�)H��8�J)�**�\U�He9��Բ=;�,���+���	
���Ve���������MEE���UI��H%wE�����Glu��D��j}���A-G��k�v�n�~�@o���������k� �G��r�(����%�#^����2v�s���m�����#��J��?����?J�����o��?���w��?��K��#��ዿ;Rp�OO��~�k_O�$�����y��[�v��+[2Zz����Q$�D(�n�gz�D�g�o�@�`)���-���g[��rk^>>
��X�rZyn�A��>Fv���%�.��}l���y��n�����1�D����!�ʟ��oy[�������Zt��N���]�V�@ � �P����z��(:d�F��`e��G�"��-��-7�S<�@8��}<���$A���">��TZ9Tu	�O���!WnC��=/���nQEؓ�D��H�Y�;�o����ɆF�Ðz�I�Ւ�fa1"hw�봈]�$��djie��ף�iA������Ջ��1�K�gf��n<�V?�L��ڢ!��iJm�=��S��8
WӼ���H�:fh�t��S�������Ŭ[+���o���E�V&��-���k������R�jZ��jY�b��!���Ǜ8>��mɰy�g�!������gp��!cF]4\%������{�R��W�jTZ*�a�1ڍ��X�d��#�^/�z)�.�����ٿ��F}��j/�z8�3��5�OB��Q %��r-�"�C��A�cc�ӭ:D�yJ��J:�3�*����0(��C�e7���ק���%��ɼ�t}�l��[�H]�Tn ���5��>���BhS��V֤uԿb����޵��%_��{�Xe�5�����jW3��2�b��vF���uv[��֮�ߗ�W�}!'�PtN�����I��t5��_�LJQ�k{�o:ZPqP�մ�;�3�]����+�W�O��Z%��}�%}]����ݜE���"��^	��z�.;��,$Qlݸ�]�ܳ��S�'�����ﰪ�kK�ucii��%ew�@��jOXK���S�1J8 ����L�y�z����Jayyx?�vyQ�����hJ��[I���2��!斕}�N6�^����1z�m)GH��1�ڶ��&>�M�����t�1�t�9}��#F쥔���y��˥EE��9*�SSS�z?zǳu~D	¥���2-��������Ʋv��b�)���kQoDwj�|�+5����	��+�_�����S?���P�5�6�=鶴�7a�q�2�T�>��{RfR��!%�k%��>8f|ՙ��*'��
���~tB����(��/�'m�A���D��H���N��o���ɮo�+v^�{��|�:;;��y~>L�ò�N0�%.�\r%k��n��bJ$ņy��m痿9���K o�炂��������צ�
A"�|3�6^)�������wcW��?�q㍡�b����Cc�555A��߿7��-����]ep≁���J���h�d�L��Kb�a^*�Rh���BI������RJ��1,N���;��@�d��Ղo����9��܇}p��]n?�0��.]�}�I�����n^,���X����0�zO��ُ�D���1��6E�uW(��N���S?>��ƒu���W�經���LQ:9�gT��Z�#>��j	�݊�ޛ���Fy{��7t���� I��a�ϻ�p��=b�ڳ��?Y�^�lx?���/g�/�����
�3�d\쥴@I��ݮђ�z��G��$>>�q��@�@t�̩DM��4ٺ(:uÎ�Gqk��k�edo�.�n[^a����X��fDt(Xx/o^w��ɓ���N��7�l�@9;\�/�y���Ҳe���2&/��vv^ aw�W�>!��5�?r�S�:�YG�Ƃ�P�H��;�uH_:��~��棬5�շ�8�g5��޽��R�O���	�����Guiw3�w^�c0_r�����тZ_gZ���6ˀ=����`�P�(�����4�w�ȧ��>���m��b���9�'����@��W*-�9 Bi(� --��-^_�Iy-O�W��d���=����fFq�<%�F���跧m�>8�:�}"�7���x�厑����d}�4g������#2mb��u�E�@�ߙ)��߿w����0�o�B4�a9VV\Z�
�I�y�	̌�����q�/���O��$%���P>x5H�@yMc��E��@=�@;5����%"�u���q9���`��t�oN������d�u���?����W���WWW���i�2y_p>/�ճ;����n���سI.��G|,G�U��Ǜ6=��
�J��f��� ri��n�ߏ�����ۮ�m��ji0�W�W�S%3��ȡM;Sb�����7s�)�J=*�������,F1����jd_ԔOu�i8d���a�Cm�=���t5����7?\��.���C���p���H~�Wԯ_K�,�ҹg�@��5<l~���Ώ�M�nb3�@ة+d����F�%�}����r����(K�&�$f{�}4A�zR��6� �(��קy�1S�|2-TM�T�|! �H���]}L�S�_l{�U��.�޷�+`8�������ҽ�ǩ�~�������Gڡ�\�|�mxǿ�,-����o(�2�NKߥ$�$��>��7):4H���C�cU�uI@H�m�I�(�ym����K#����#��B�%�:�}�D:���L֞���������O�h��/��@��~�;�Sjfk�-9�j}��g/�å�^ȵn���7�7����ȧ�d�ͩGդl��ݛ�5��Wu����i�s�~�y���Q�����Li�
[��Wr���!v���=�3A�G�KW�uN"������T�U�h���x�u)l���/p(u�BV郞N�3�M�|��}647׈�;��1J��{�����ރ��5Q,tǞJD"d~�!A�s�2y��]�*v09jd��a%��Y������nƄ��G�MK�:I�+@���+|�����V�V�����3$zqr�g��j~�Ϛ��j"u�G�i%y���:?���+�=a¶Q^���D��6^�#ؘ���6��L���X�V|dX�=�~{��������������T�yV��]cƔ��)Jz��RD�]CF��f��>��>F+�~E�x�}��X�6���>�W���S��g(1ѥ��'�^���_2�N�F���zB���ꦮ�W �Lb��ڶ#���_��~L���{�*{�oI'�J2��H����3�cP>c�[C����sMuc������K-��];�cn]�*F��u�#�(?�W�hJ���s�5�����]r��!EҰ9Lf��v�BI/"�l@i��lm[$wj��|v�H��}�y��NM�������?Np~�s�ԩ�"��v�/6�:u����sp��7�����v�렑��-�b�����"<];��u�k�%��6�����a#�A�X֣�]���u�9io������Ա]o�/X��n�Z#}�x���O�"��9 ��7��:j���]��v�h�HRN����x�5����/~m�z�T��Sj�Gc�˟߾}+���c.�q�$�I����ڷ�`�aܩP���0v�и��Z�g���P���N��������^�J���'v��.��AR��I��5��.�������q��Dۉ�Wg�I���͞ﾁ~~?҃��;-L3('�?��ڽq��#����A��h�'o�T�Ȳ��,�?�[��1�}j� 3��lh�fi�d��D��K�ס��x���/�)��8�:�2A71��l���~�T�X��mW �h~��r��&+�������
vRw��%�r+E��}����",�C��~�n���������pq��U/����.Ɣ��<���;//���q��RPo�3w[zM)�e%�u���*�O=�	���/K�P�xdé\R\�E�>������I��=�R��z����,???1�������.5V�N�������:�z��/N\�U�Vz��+���x4�^�(��j�gUv;��1!e�{Y��q�	{!Ғ���ޫ�d���)�+'�\�;`��٪ը�s�#^_b�}i���ig���Cx�B�A��8��T�dc<]4+���Oq�A|{��,U�Ђ�\<���|g��E�%�I%S�s4���e��'�o=̼�*[��̱	q��/E�W�b�C�;����O�gd��G�Cv�Q���_��*�k�w��p��zW�p��5t1+��{��������XBO�-����f���>�>mTv�Q���u��%�rT�)�̉���X:�J��ly`p0�؂|�ׅ��-�v?���ॗ'���P=��[Z��?z���L���I1a��P�L�W����%��;k�.��vɘ�km�y�̘�f��D�`�PI�8����L;�d}8��Bgl����B���Ç���mi��'�+�jl�=Y�<%YՔ@�
��N���6_�a1����i����h��»w�ʁr|E�z�a��.��>]H"%�r
��/�Z>A0�fc�pЉK�3n�V�x��]1&̋;O������W��le���̩����09~B�xo����d�BӦj=B|ٴ��h�����������-��7-��'��P�����~��{�r->12�φ:�X_��o��"׌���]v��)5J�)ux�l��w�21z�K�l|�um�1���ظ�i����Ȉ��J��l�%
;���0���;"nW���ߒ̄!<���}y�d$1�����VV�R��lL}�B��5�h�ue����~7m�%4i [�-,����p��<&�N���VZX��y(Lhw kBBuB|P� =��Iz���n=Ո2oB����4W%K��/3�����>�'�Vr�sh���Y���)�	��'��-��?�� �W�!#���ɶ Sՠ����)�U��:�]д9�����=���؀�����vn�^��9Dx���7���BB�ڞe�W�N��y4��̹��k����ªgb����#`3p���+�����$�q!f::�X�����q�tҍ��B��zݫ�Ay����T�tL
��UnA�h1eϙ�Y=��qHoR������zi�t.��F��QI��e���o���_ٮh��XS��� �5����U'hS�q7o�pH|�jŧ`E��>5U.��S���d�=�\0\P��5�x{W~�k��ff�1*�EW;.����I�z,%��P-.��*�<�2�	f�~��s�&:v9۾��{��L% | ����DC�ԦNiN.V�5/n[$���'Ga1��\�Tܛ��K64R$s�� j���<
3J��������d6�bZeڋ�ԟ~������W��]�Q�X��-�1���V�s$L��ε3�@]��
y���-���dZf�~^�#A<N���Ҷ��o��K�B�y��u3d�Qʥ���t���x��?F�Μ����L�&~����k��� @9݉v~�� �&�܍W���:U��j�ԯ�y�G��x'�Ԧ٥DT,�,É1�A���,�裢Ymv)Gݫ���l��?S�/��Jx�=���+��u�������������R33��9�v60����\�|�Zܪ��-����T���9k�ݕ���j�(+iY
��7w�^�1yP�p�K���2EO�p�L6��&+�	�t�e�[XL��Bo��h�-�?Wgj���w<t��̭�%��|�&���W{��J!����O?ohjz��b9P2��
�<�X$�sR�|D����"� 5���&�ZA�����/\�E%V8ϾL!�V��EM^U�t��R�Շ�G�=��ם(Ϻ�IS�z�Ņ- ��"9��X)���O90&�]ߤ����Q����]���i/�����߾���%���z5�`�������ut�|]����&�j�|�2���	kn �cINy����~�ւ�h���������G�Qd �U�@#�ߎdZ�Ё�QTf)��
\)=|�Ik��?�f��x_��@���}ݭ���)���wשΐ?��/@�r��X��wH�)��w�G0.=K��}��&��'˂��|	�j!�JrI��D��$#m�e�t��;��4M�L����R0<�o��,�N���9�ã���AV�[G�v�қ�NQ�����WZ,���龀�t��ڻF|�:�,�;�@���g��>�ͧ�\�K�B�݊��B����w�el^IęcĻ�a�%Zv�l(dFT��7�$YE	ֺJ��s��D�u��!�����C]2��b}�|���AX��᪪�;T"O3c
v�@��{&�&��N�/��s��ښh��#H`tc��Z���ZPo9�8�+��6��iأ������rǱ���Z|{{� C�%Y��.�w�UZe��������}s=)����v��f���dE��N�Āu	n�&��r������j�X8(V;�P`�E��< M����s�eSS��[&x�׸$�^����vxLte�	 ۃ�YZ���[m�U�	6��ص�x^�10�v����#q':v��K�1a���L���C�gW5������΄����J�V[���Z?H8	�����=9@�q�?ؼνW��~T�8�F8T�KŲ���j�~��p��iְ�\���zg����h�ג��1�rM��gP~��ОK�Nz�$�;�o@��{�<88�����r+�C�Y�'�e3�A�� �v:�P$yi�}�
��p�j��Ǟg��dvi�� b�A�zT׽�|��1G9m� �І
h
R��͈�oO�`��HO�8�K���vh
�╘����8|Ʉiύ��'[-�_Y9�]f �{z�����Hp��m��� X^U�R$�X3�u;}��׆q��o9
����ԥ13$�9�iH��������*�	��$���t���F�qH	�P�~B~6Izݙ���z.����&?2I����^3��pO����WV�(���c2&#;�r7�#~��3):�k{K�
��g���u$��Y�Km��˃m��]��0:�� ���0c �����Ԝ�z���#s�&\x9�?��@C ��
|�ٲ6���#����8iZ�g�G}
��>?�ӟ��v)4��i�D7�	��a%��Ɂ�"أ5�?�	4�bfDؙ�&&0���Dػ|P�K{!h��S
�9����\���������0��Jmo\*���B���*��A��N��Ć��3�=s�D�t�ĉA}F��φ�p�/%�"�J�N�I�au�~>>>�(���60G8Qw�z{�
�� �@�UE��;$�I�Hh�q �W|�ǝH�R˯ܭ��Z���k`��1d$޻�L���KM�w��� ='��g��w����?��o��r��3���R�o�3�j�]NhV递�U�����#�$x��p[���q�/�ʈ�d!���z:H8�3*/�#��M���HH�)�����A+�Y�	�@"���Nr��[��V@���H����R~���HY��b�L�����EY�M�` "A o8�R��-D騯_Ǵ����}�R�Av@����&�%���Ll�WO�4����6$KDt�``p?��#��z+�3�0e���G��u�nG���@���/!Pf��u�Ig�\�+V�4�����@*�4�0p��P6���Q�c�4'h�l(�C�]ZҪ��4�%�����3��D�ZD�"G�9�$(1�Z�hH�sC�	&���i����K�xo�CZ���`<Ru�JRo��9Нa¶����EB�*��n[��,}��q�����o�$"�x�Xm��OY�Xxe���`.�)��?4��E$~�B�h�=xm#��?��Ř�×SnwWlד5�^˫�c(Tj���R�.�dh��0{lҮ�r	�:��Q��E�I:N�c+�P�J������I��,5�\4���\e�Q���'w�K?���g���9�UJPOnY	8t��;t�#�c��K��F�9h�"���o���<fP*���qa��������u�)�M�d�R�����|����C�k�%����Z���o�a8�4Ĺ]����Z�D�A��_{i�V˲�YeglllE�������*�4Ǌ^L�g�Ԧ�+zpE�WW�/�C����>��(5/��!m���mM�\��D4���|��u���::�F0��-�So��.M��qS��q�^vv������΁�@{�S����OO�ó�Gq��k!G����L�j#0�${���~5�w��ݑ	�H1��[�����ڨ8��vcc�wjjʠ��1�rGVv*��>�.�Z�3k�bc-Ѳd����=�O��<�k����lJ�C�
��G�<�ۙhI�<;u��B�Ը���$�ѓʢ��<EX&1m>mD�=�iw��iY���F׷�����#6I:�x�$
ŀr(�lX_��sYVr��6��l1�M����!��s)��SO>�;���.34�mB��sŽ��0�L����YhVp��k�,��O	�R����˃��r.̡S�X�o����.KE9��x�y�x�iYs*�|<&�
qb��#�~/;j�������~�Ӄ��Z��;b���ٹ���8����y��!u��8G�P�WV��i�����?�Fa��%drQě���!��if&����=�ư�).&6����w��"�Duau�0�8���'��>�_�B�dm9}�K���ѳ�a?�wNݘ=�<���j�������f��jY���zT*էǽjS�1�3�p�����vò�^M�1(4г&σ�

>��LmC�[�d�����;�e�Ч���);N"� �m���VaՋ�j�	W��������BƠ���"�A� t�`H��!���0D5�n܄��� #����G�����s# ��[BU�����j���iG�{��D��v���ުA����+8��;ՙ@U��M��N�~�J�Z�Ri'���cCx��Cehg9�F�ö��Bu���c�}�i�[��+�@�}� ������-_���5�ꓕ��8itQ�Ӌ7���R��z��' S9�����Z�Ipyy�܉�O���ٲ�a���,v�J���]�����r�\1
��Uva�5D�̀���W��i��p�Es�J�^��5�ɼ$z��y�2ys���Y�g�ѢW遉ZN	]����i�� +����X�oՔ��}����ҁ��]O;U�Yx��eu�thЗ�c���2|�N� q�+�����Z�r��yyy]���p�B�~�K�H��I43X��u�R_T�k��������������g�	��
���*�F��������D�׋�"�8�Qƨx�T�ewo���{ٽ1��e�4C@��'l�XX������&a� 4`�w:R�!��l/$�~��A��?
5\ ��C9���_�ʛ��K�Zp��160Q2$���1��"�**���."��D�q�h��.�B�b��#a��s0�J�ZO!���g�c%�H�A0�Vk�+�oT�=O��x"�u���ɩ|����G�����bյ&0���V���g��H- ���.̃�O���6�7��臬�LG��~_�nUs�&��	5�&��7�~.��ŻQ���-!�yb8`3
�G��
��Uh��:��?�h*}��^��N�f���^��̹�ϭ?9��W���@EO��1
ȡ@�8;���Sz�^V���HX��.--��_,�j�3��`:	b�9�S~�x���mgc�!b�W:(���=؎��ph��B8��I�-�����D~�0�p[CqQ�1]�U�������r�mF�+1~�����)8�}��!�� D�µ!�פּ��C�����i��l���b0�ap8/d���;�&T-$�0��+��k�"&x� S[W��Q �-߿_���ǃ9k�s�aп�n/����� �����C��0mK@�s`����m�{� (_�a��*��jȩ�qo0[��tX���\V�Y��qbY䶶z�9pBW��8�� ����8�@	m/����/l4#j###4bḋՋy��]��S�����z ��UUU�@��sS��ќZ ����R��"=<�P�g�Jw��3D����5S�r��1 ��҂�9Й����j	{�����?�Տ�%noo�g�L�:#�$`EcJ��%:�� ���)��?�mi��xx�� ��I��m��=X]���gi��2-�*�K�9�� ����5@(��@�=�f�>|p��R���Ш8��Ì��EC���?(I#p~��Y|D�����n�n8q��ג�YeIz��#��I5�e3,��<cKkd�[qя�4�c�ʢ%���o��������c�����u��т��j�C�d�h�'���D�ƒ��$N����+8�_�h}�ala�ejjj�\KM}@�xV�RB���y0��]�����3�綴�ݠ;Ȑ�:
bN2��T��T�l�A�>3�k�]p�Mh���(*���RV�g�3��Vf_udd�g�W/���l' Y2��{)UW�R���K�9-�����a�櫓�?5�_8Z�����u#d�D�)�얓�>� `V0;ڒ]a ���f}�6��x\ڞ�lS���KD�"	�Ԋb鱢����"6�S+Ɲ�8:?�gLd ���"�[��,�����C&�U,�jS�)�3䲬�"�KcQ�Ȉ,� ƽs:�pzv�����u��5"�ו�-K]�ago��Ej$����'�)՘����vq^�\Zy����P��F��P�����*B��m�98�5_v�� ��\U?����PkK�d�-f�L��Q�Ǉŋ0[�W��D�ɢh6`6���h�RsQ�vĞ��U�J9݌��}'�6�H�c|FƩ����QY&�����JB�KDS'�>_>.�fZ�^I�}�S�~QC�2	���"�$�� $��'�����,J��0<�vʛ�zS�:����y�O�m �8='pG�q.M�x���j%��Y�-�Ɇ�/_�v�L��魹{x���l��ԉ �@|Βl��şȔ���2y3�C1}?=����=�^�_����ء�R?ڱ.�Z�K���.��Ʃ_�K�*�`���B���!��xaBݶ �ȃ�����
B�z��w�0�������I>����60���x��]۩�1 �DB��I��/nG�Oznm`uh��Q��]/h�5�/\����]1>?h����D�B�AV��f�~������v1�:�j��ę,A{�_�s�6'��d�������^R�0grY�	�6���l(�mWH>-#^Uh�pN��y�૜��5������[Yi�(^=���4z�I������J�d�"��"�J��ﭵ�ŗ%���%�)��vgd.9�!:��,�whIWw/��| �%[��&~��9����IURg8o�������/2��T��>��8��g(�������|3�~{���1!Ҍ�]��E�����X���/��y�����i#>��ۙC�ƍ3�r��V%5N���}^`�~y>�걄w��|�ݶ;�?懬\�ϟ?[�\,l_��V���v��+� =)�o�m�p�L�ً�b��bi����������C���A��?l�Ҏ(fk�ͱ��g.����������o��NN��H/4���w&�»�9d�A	�ss@Lk�. ��o�*%��Ֆ�hyc|*����N� ��V}vw,��8X����4,�>}ڊ�I3�@;*a����;~����$���Ѻ_;~%���|>�B�0����Q�k�ĬIy���TU/YN_�qP�y-1�qWup0���~�|c����o�z'���]!��bg[88`�H����BX@t���-[�EmEE��O_,�>��"Q��$�l�u�O>M;��9��;��x��3��P�%�;<��$ǯ�.�ғ�h��T���x%�T�j���\ӝe'�}E��-/��&�wW��`d�.h/��Mkoo�L3V�+��v���jrV��
��Z����3좳��5{��:Ӿ��-��	����6��m�����>mUTo��ƪ�7��Ȉ�#C�)�Τ�6�v�����ii�cCC���#�/,�D��2�x��;�q��G#0�	*�+��d3#t�����u���`qn×.���:T��X���xy��������y������3V�}�K��O�=�(�����Z��̣1��1�]�	ݭa/����Qx`0�ѝ��'_��DJ�^������{�� 
�oS�o������j�O5�E��#X�b1�w3�����<��8�(c�/×�u]��Ô���j��8�I�KEVгN�/��[\�9��4����o��Go�}����{��d�Tk08J�_�)l���t%�0w1���AW�\����h��CJyY�t�nD1��(��ő��u�2�P���<(�Vm�U	�4��i�)I:��]䕶4a&p^���/V*ό��[�m��5�m���-����\���Y�����8Tv0,^��(��%�,���Py.\)nWTbtw*�Q��D^�c���o	��*a�B�-r2��B5U��,���H�����/+n��h|�����8����bK�Ս~f9��|!y#��-���p��]��n�u���W�(:��G|R�Ҵ��t@]C~�Q������}cn�<t3� ,��������J�'��y^:���h*�e�d:4�r�<��ۭj�f��%�����z^/�p@pV��}h[M��v$ȻAtNW@�{�B�P��ʣ��Nje�a��gW8��|�P�z�@4�*�2�:�ٲꐢ�zh)m#�z<M{z�s~~>��"G�/�t����{gf��&��>{1���i�Ho�n�a:U��n1��2���MN�K��g�yLB�����E�k�[����FT,��.X�X�EƯy�P��g��B�^̂�&YK���"���ޞ�7zEmkk+*:5��K��v7B�-���ކ�t�w�h��e��h)�Sq�m7�^�a$�YV-<oZ	�r�L�nQ+��;�}����*�:ݣW��|娰~_3�_"���Ғ�H�sm�לU�!d��(�ﺖ~u�ӷ�k/>�	!F�K�lpQ�d��z@M����^T<R<1����|��XY���C_�_^�Z�r𞥴	���+�G/��u����G���T�����$�n��p�b�4,S���@yA�~�m�L�{fm!�dv�_��nxf�����V�JT!0��
i�X����{gE�]�!�B7y!H���]|KJK�4C/�'m��Ϫ>�iG�:�_㿊��Ċ����30uu�W��˦z�e<�E��7,�L^sꋸ�����]�M�d�;�M����m{h3=*sɼ)�(�r�(uq��v��Z��c� ���w�'�uh��[[��Vu��_?E��W���7nu�՛�~��(B"�$x�n�퍞}ɝ)�6�<���=�C�I
�}�T;�K��_�.�	��x��*����__��Q�/�O	I~����̧u�]D�����+cZ~?1??rَ��6Gi�m`��UW7�vX^M���0	5Ŵ�~�^����;����Qm�ů�5���E.N8�N�|��y�j>M�fbu[N6VV���ݚcag�R��!��]��۞�j���㳢vs�brrR�![�i�>H܏�T��G���"''L���2'^����=e9Thc��`(�y��Pl~y-Ă���#H�K�|{u��M���xUU����<��W�Z�q3�b�үm��J�|�\o�y�j���(浮��_�\g�V�HWY󈦣k

��7�_�9r�-��̑�,	��#p��q���40��M��e�r�T��t��)��D��9�I&���8C�0�d��$�r�a\tL-k���I���@sU��A�)%�e��GJf6��X~^��`���77[ׅ�A
h�k�U$ڎ}�Mx���İ�*oP^�fF'���'�GF~��И�4:�p�3]�I��0�B�ZGDB���f��Tc�
<��"�C,�����J�x���B���&�b���ԓ����ya�w����YSNmIwp�|�����	�П��۾�����Ť��u��7�	Rv�ǹf�т�Ze�Dܕ�������G�a�lQizx]����g��v��&�ʲ��-�bV{�m;h�/'�y��������*!s�y�O�?qp���9�-�fP��$e,�TzT����$�M??�W"f�>��R��۷�oyg/�l-Z*��������$S���_�����m���5�J����b�8����Hg_��Z�7��{�R�ق��U��M;zN���Ɵ�GEF�p<�LED��G�ٟW$8	�w�/<n�8CnEV�g}���ʊ���|�Tu�p�gY�JgQ�UE���uW-��J��ɷ2�J���v��l嶜��,2��@��Ϗ\�R���`MK���P����&R1�(�d�2��!e�W�p�T�����<
���A飃E�����%�[�4�	��Y�����_2����������͚�^QS!_J��gN�=�Q ���ߔ(ͲqdTϲ1�f"����M���d�kꌋ�M�1Va�����}]ڮ�����7'�2I4�?�r��ツ��;]#�;)������{N� ��4.O��"A蒳��HUެ��iP}O������^:v<N�]��V�����t����#���M�j�(*j�]8xIA6�?���P35�w���J W�{6���N��`ͻ���3͋�@�����#Vφ�8M�Ύ�ݝ��Ⓦs_Ę�Y�a0v�J�F�;� �5Uՠ� ���W�yłI���tcc�A�d�hM��-��Ԍ4�x)��⵹K6�eW?x;3�-M���D :(����3Cg�~7�~��kG�_I�D��}5�E��س�Tk9���~tc3\���.���ʯ�<�+~t���AAa5�������R���Ϟ=���;Ӧ4[sӨ%�z{�����w/fV|�y5��"c��I���O�V�|���o�^���;6���%ݎ��LҦ���`����kN����:ng'$$�7.�-b��!���[
����D��"f

A?�U��>ǆ����捏��O&�5��޷m��|羳��_U59�0[�#����}��	��pI�ҁ�)N�'�Ș����eO��J~��a®���-_g�8&���Տ��SS�0i���ϧi ����&�����V����{��ZrC�G����3Z� ��v_�ueKչ�b�w��"l�YMM��L��*���LG��9��}�2<Q�_�h4��%j`@5MK(��Z^^N-�5S�m�+c�Z[[�����'|ttt��Gs���;�a&_W��T��4�a��-������¹�<�$��D�����*��;�MĂ��:]�s��	�����}^I^���Fkk}��2��m�r�r�C%�/S3ܳ/C�K��h�LnRǍ���R���LO��;Ny5�]7S��V׺�>N��nG�Ly~ֵ��{��w|�c�I�l_)�̯b;��������B� �讂���H�N^��b�w863S�%�UIz~>t{�7]-�~s�f ��í��=�Ǯ3���*�7?��.�pޤ�d�Ͻ#R�|��	�	 L�ϴbD'X�xC�SL�mVf빲"�f]����D+��]��`&$���}���Q���m�o��DD7��X�stt�O�W�[�pG`4�W��Jf����ڌ�8������ny�^Ϧv�Ì�n�g���۔4��G�V;8�W�D���j^EO\y�ak��G�Et^$֊�5R�@U���5R�55@�f�f�7�%s#��Ri�G��:涷�VZ�Ö�6�\u�%δ/s1k�T�Nj^��ˣFl�sj�Z�X�.�D��	_|�]�=M̖m�ɜb��ɔ�o�O�d��bĠ��MV#���lx��0��ix��;lmL����G�-�Ҋ������ӄS����q���gς�����ȸ�m���p	jVtں�ʺ���$�����yz��������P�mۖ�$�B��Kdk��J����d�!�`,3��Ȓ��I�lC�!�w��`��/��X��^������s�������w;��{��y�W]W����*l}��6��ዽ�"*而���a�Ηp�y��o�=Vϒ�5c�uAd'o����'�|�����(�Y�u�����1��:\][ە���h%5&��iXx��ׯ�̓Y3�xTw���o����K>$XzZ:V�{'�[����a�-���%o��̱A��fM�P���Qߑ��*Ć����NLOK�Q�)�t�T��ST4ڟ� LKK������~���4��ĩ�s�A���_�/"�R�O>�N 
�/�s����w�N�测��ivuyGt�;�����I��N����K�_��IK������������а_-@�	1��[u]x�F,��eA��H��d����r֎upI]�cq�`��_�?{B-���� ��_FW����@_vht�5P#�,��d�[d��/W�O��Dβ������frA9���~*��RΧo|�I�'7nP�f�;�����]n}۽ǟ����{"�����15UA�G�d]piXA��۴^��y�0����Q�����!T��ړ�&��V;��֭@`
ީև�\ ��q��7�l9o�j|�k�u�r�x1�eg�r	�T�̫jv�+���ٜAs�ȼ��{u�Y�56��+�999����ccc�y:��K�o貊�A���.�"I�X]�Q�;%

�>�>*
�^:M�.�6W����VW�ҕ�փu'�y�"��?~��CTR��g�h��)�3�I�,g+�||6:\���4�@ T(D�421����� �Ys+�b�x��E�s�d��c�<�:����p}��ę��ɗ.�u��֛�#{GnO��a�O�Ji&lF��n���3>��-��Г� ����$�<�vP�?m	?-�,�	
-���_��}����Z �v��+,"�g��@ۘ����!
�sriǖ���wv�RS�n�UV
�����ݗ�'�zPe�BK0	�Wr�F꣦�L���<��f�Rp�����!U���\�gRKǞ��ǻ��^O�2%f/��K-�lV�l��s��
= d.d6T=���?N_��75�{�]�)�/���R���pR]~k���H��3�!����Q�N�Ka����_
�[}"e�^����кZ�FS���.pv�Fw8:J���nɨ�l@}����#7��{�1���3V�M�by�����:߅���i�t/�wpA����������ֵ	��:m�L�kƉ��Ju���9��q?�ZO����[u���S�^���͒��0u�M��!o�A�i��B&�8v����U���� �����AB���lC������s������Z78]A���#����觍�8�4�"تX�"#�F�^��
O�N���q��*�ݍ�V�z�w�+��M�6C�^������o��0����T&���O7z�q@���ܺ�
}t�C�>W���l�P=��E���p�{L�p���k�y��NL���%Yk[�p�
_va5�oA�`{���;���D�a];����R:�߿m���l�����]G;�E^���RZ#;��m+�Q�≲0��ہ%�,i�՚I�}Ǻ����sH�����8�-eQ�ǭY xH��V0Ǥ!���j�}�� ��פԵ��}E\��vG�cΉ�j�PQ��,<钅��ڪ���g���@�z�̳��C:I"��T}O_ߛ"䠳�������pщ���LNXN�r�鯁CX{��ǣY���J hL��M��t ���u�׀�����v�1�VdP��u*M4�Z�DIq0\������}�&�#�������3����}W۫z�ʒ��e翓��:�Nobٺ��M��#I���Q���-��Q�����	�e���.�Lh�։�AGF8⠁Ï�̀.�%��3Ï�����W����V_KiK0ƀ���֠���p\�n}��lA���YuLr�j.2��_[��n�J;�LG<%�������}����!@�GEB�:暶�Y>�ϗ��DT$A��� ᤯��9��1Ѻ8}�b���X����칬���@��o&�H=!�|5��m�C	؄�@�;��̧4���R������:��x�o|�(��q�=O3��L1��ZK�K�>��g%%������_ߎ�u#�H�̷�^��1�ő	j��^-F���9-��y�;fbE��"X�D)s;�[����'+P���(D&�Ԋ6��j*mu�A��ӡД��d�|�/G��TA��ܸ�"����v�I+]6����T�C�}6��n�j��`z:[8#�N4K�Q���k�#��{�cʳW�G�}��C6s;��~�\KS��J�K�_=_�cM���lH�������u:�~��O�d@=r��-cԑ�	���t��U2�v���A�}-��4���@�e*l��^�?.��A�0`1���}І�ǋ� �]n2���BL���y�|2��&����:��%��]\;,T�T�������{򽛋���Yp:�a�h�IH(c���XO��1ATU�e
*�Vs�0�
�ЇYxI�l��c�b��%��T�hpW��̔��-��nZi�
)_M�ș�V�%�VL�q��[﹒��-�k˯��#JTɘ�A�jʇ��	ÃO`��� ��'#6}�f@+S��1O��ї~I�w>��9�B,ֆ���U/ٿ�{���RC89p�;{g��7e��X.�'�|�r���AN��NB�g���44��^p{c��hAN�0�ܲO�+�*��C��m�S�x�I�m-�u�c7+t��~Fx�!�\�T�8��W䬀���
'��j�P@���j�V�C�Dj�W�U�R,Z�L�JI��ED���\"Q�5*�JZ95���5$�
��FZj�0�A�TH��&�:`7��,�?��'�>s�8<�j�Y_7uΑ�0?u�N`dM��޴��)�ko��ym�Ul�̝B��Ѐʵ��i��k�E�X'��7���n��+O����Z�f�YzIv�{mk���hA��1��N��0���Y���S�y<8�!y��i2�l�#��6�:�ף�O�g.t��l@�G/T�3�����|)�=Q�^�_~����Z6�[E*<�����T�k�h���hDk(L?鼳��QR�J�+1��yHObaK <��5-;}�ߟ��!mf-`���
�0��S>,�MnMN�{R�Y-����y���z8��K!O�H��ɻ�nV�ū�/�xޚ�ټ��5�Q���ثP9�n~p0�K���%�Sk`(l'I�f���d�����������\�ҍ���5���S��K�3t�w���=;;�BF6��Ê�Yi.��NN�/��R��L"��t����z�V������]'T�������G�dA�*7�6޽�#�w{���Ҩ\_�&�W��)h�y��r�S�t�{���]t�8wW��|=~n����ByX�l>��6��[f��Ӷ�/�f��ш���>CͿ�I�p k�c�1o&��״-�����V�Э��m�WA���~1w�h�n]���rw�V 3�l
ݪ���e�.��{���E�����8&_��˄.wa�T�� n�I�?�г���\� �Kg�ZUŋF�b�vƼ'`?��c�%EV��RHp3*b�@��h�lɫ���ڿ Ip���dz��rj����3O��o/KK�ҁ\l<ǿQ�0d��ȣ�;���	p5��T��x�?�JR�ѭv�JC�~�)F`N�+��_j_}��xBEYjRG$~/}[�J�E�r��`l��؆������c�4 K��� ^L%���X���]/��Cs�-�g����K�;���pn���~^eU�����d㗸���'y�;�%���W�TǤ��j`��	�[��`�7�b� G4��X5�y�EH���	�x�SM�DS7ŷ�L�	�ch�{���m����^�"B�ǁ��	ZȂ�iB(�?�X�[� �1镜4�l_�w�w%_ce-�6r�'u�
[����YK|6��xx�+J~�<��3���&{{�����p�W��-��Ϩ|&z��Z�hmW��,�<����)�y�8��\���Q�UY�H�9�Luw{AN�҉g`����MD�t]������,O�3�����XDm9���_��s[
����:�PmU�Uk�k�Tqu��먧є��)���f`�Ͷ"+�;繧wC(���~�/*��}]����K����_���|l#�5<\.���L���\sHن�,Vh��J�:?���\�ΒcH	�d����v��_���v�ԯ'��ٳ��8�SKu�۸;A�)�	#.��{��[�v�e���A@���F�*�>��ڸ�Ɇ:��7�:"WR�~�g_�	���ʉ�����&��� d��wv���+���x�2�M*�1P|	�G��@}jR��T~9D��@zꍐ$�7s���W�!(b#b�$Z��%?P�![��'n	�p�ygΞ�F�w�~%a�!RaO��㙙�V��NBS/U�@�Ƃ���aV�(Km5:<��M��T�iu���2 e�9����(r�Gϩlo�@t�=��-�z4�ǳ��'��nݶ"4�RZ �$o��pcs�$��+����zo}���|���^9�CLK�-�hp�<�ק��L\��	���j�9�o�X� �=kvf,	���������/���.�k�=���p��\Ǚ����j8quPsUc�&��ZˍN��������=e>9m�aoݖ)[ZN���O~��%WE����&��NPfk��;�y��A��s_?�vB��zd����&��4����9���pU')NM��p$f_��Ƕӆ=9��dLB�u��͝�^��i��\p$��'+���.�ؐ-;�a�����톙	k��
�zd���gl� ���M?�K��Q*@J%v��D��:���yX�Ե��6��j�4õ��_-q�f�z�t0���eCu0��Q�T��/t��ƹ�����U�2�����Wj�t����1������_&����@���1�2x�w������;�i���9�}�1�g��ATm��le5�t:��D��_?��!�|�r�J4T��^�������`�͔���8H摫�m�7 {!�|R�뀲C�	XO�MIt0~��l����G;Zs��`��BsL���8�EG���MO�1��CO��%S����%�3�7��w��>��{?�=Gb�E��3�BiGNi5/=-�*z'>����oxk���a�ٹwb�2"nVSBΧM��'i�ۘc�6i��\�ޒ��)=��z3����6����]{Q���?d���]��x�j9h�]E�\�eZ�k%:<��D�R�|�X���ɴT?	�+�-��t�|���Gh3��j&{Xݠ�z�Ò��`|˙\Kg���r/GkH�sV���P��>W�P��M�zx����&R��
�^F=�S���'�����0��}Ү+ �VR(�Z@vCS��Q����x��L�ũ��e�0O�5��/ �e�4�ڋ��㈒U�U�bU�}�7�{��F�S������!�ЌH�!0�\�a��|�<J�Fw�QUZ����s��q�of��%4�}7:V��j�==��rc,7�,�$yO����L �*'��<��
~�c���x�o����Q�����N茅_b���:��u�ZA F�]B��@��4Y����	T�N��ǉ��=�{���e����팔N��C�9&7�,��I�B�HWp5�B����!��aM�28њ�
��F߽��;���ǚ�Z� I�� �����Q!sۻ�o�ps̮e�*<4ѰQ�rW�m=�;ƾk2�+������)��G-z�_�,���[{Rv�\���*Y0Ki��?�s�yz� �z_��IW+=<�t���Ljj���y�L��<�v�稽�e�q�+0e��jc dq$�C��j�}�F0�kD��F��\�����F+O0�����a�-X)�Մc����/� �����p��NU�D�4�t���%���{�ѝBUa�D+��k��ݛ�^��j��0rȤ�}�lр�w���p2eI��U
��j��߀��Ig�u���s�N�u�i�~-@G8ID�7	�~���4d���`���5���1�Pؿ��H5����U���FA(�W��}��|z�3qϴ���j+�l�F���}潙�n��S��ރoE�,�9�Rޘ�9��i�[�0�UU�%�ێ߇2g $�@�i��i���˞�LN���kq�-4oDEy%
M�x��ޘ��.�O�WzFfG����,��v!_���^#̆�	Ke���o����Rz��8�5ǽ�)��uz܁F��^�M\�����.FӠbA98�
�+(�$;�j"L�tv�G7�zp{�Ѱ=W�u��lR ��ŽV��=`^�1đ^��1�C���W�\������b�Z�7{5�#���
�?ծ��ӆ��Xߵ������_\R�J=�GF�\��U��ʳX���B��aDnw�����9��ȅIa��f���'pO;ݖ��ﲲ���j�r�NbJ/~��Ef�_�F������ʬ�~m�̟^��p2J�JY� D7��_��r_7�yS�c��V��y�&)�����~�ђѫo�q�\�$�����HZ~��Mo��Z���p��o�PQ]X��`'�B�jA*0Fd<'�!�����O��pb�C昔c���9��/�h@�n�<7てjC��߃�QIv�fn�e��U���tt��x����֮���6zP���D�����ϑ�ФLd���`i��"i*`b�#,X����V�l�T2�/����.b|�I@��I�W�i��D6�b��т2�N��&���ݕ^ln\�:m����~trI���L���yN�{^=�T�(F�j�b�g� i�6��dӨ���qK[qo�@.��oS�)��)e�:o{��U����؆uҶ)�jL�̈́��#~�tr�Vߌ�a�E@� ���C��Wt���f]J��
������u�|c���	�3+�^�/An�}�7���E���C��?���Y;L�ʹ5��J���~+�k��Mv=7q`�v	69z�έ[F�	���:3����ϛ�i�����Q%M�C�E��Y΂��gFۋ�ceIΞt ^��_?�r�ɹԻWՔ�"z�V��i;&�N�6��:�96�T��5	�s��y{	�j��R�Z�P[��b�\�Um����yxb;�R�sCA����z2� ��V�J�H�~�fʯ9z�*Z�߆�44n�Z�JO��twTF���G�ir&��u3�UG��C��`"�'�x�z[��#�.	�R���c�49�튠���P��C�,��d3����ՒY8Sʏ��W��"@��}}ө˙AvJ%����fΖۿ[����Z���OU���K��}�P,��f���ԡl�es�ˮ��r�z�8S�؈�����-�<,?4,�\x�U�Q}�	���~�zx(
|�*1'0o�=��- ����xn��ܤϣ~Cy�z�`�>�N�g^&���� rl�:����\�!�)��"m�E��5����J�/ub�`����:���1�����(�Z-��״bҴ�VTM)�I�>X%�T�~bU,.^���K�����t�)�̱���
L���-;�r�X����rW�酇�*q�&��.�{ׄE�b�h'�*rS��#N�.��T��+���O�jI$R�-�Mbd���
��u]�Wo�T,�<���M�aI:�ՠY����<�H���t�o�;x/zo�Hl.'���a�V�e�jK�z7D��I����u���V+6�9�����3Pi^AZ�>>�Ws��Kp�G����1kt7��XD�j��;��� <���A"E����|+	�]XΌ&���%����{ɪ��aۏI�!�`V�@��Y�1[@f��$Pe�:�X ��cÏ��ӳ���y����u�~���v�S���Q���E�t�ܛ!��]�7�Ee�#-�D�T>�&t��yǼF:���UE�U��&X�%�%��aU "�m��ľ�#���r�r5�Ӊd߭�xڧ&F�12�Ò8��~�����hGaUz�5�i�Xr����fi�P�ͽcef9�J�;��l����ü�Wac�ל� �f����ٕ�/t8o1eS��E�u4vW�A�XT5�
��L��A���ϒ�N�
�];n�-�h�7{�*��˙}�jb����U����5V�U�B˟����S�O�Uu�
F賂x�ӡ�X(R�(�� 6zh���s���t��4>5k�
�p��ܹ�B�����=_]u��� -oT��v,����G�6�s��������6��"���
�C�ͩ3���\oE����~�ȼ}О��P�k�b�m�!�0����kc��*�܉
�m�FM�����$)�{"?iiE�qau䯚�}#���3���������knש�
\N���T 냲�.8�B�ە�_�Q�A���5�D����c�ĶY\a��������^�����O�iu��@K�4�h2��H&�j#��V����P��F����w�1����s$� �z�,�:��C��x��w#W=����L���=5�֐�~�z��"�5V�J�.�͒�p���.;Y�������[|�c���
V�Z���T�h�]45d*�z^���o�x�7@��0�?�)��^C�͜�;�kRS��:/0�W���;��Բ��U�VGX�������8�u|���0�}�~��?8��ƺ����un������k}p]So��91 ���C��*������o�����y��Z'�����ڽ�U7�vc��҅�rp�eڏ* ��e7Tԏ�!�Moi���Ubo,�c�@��v�G��de�뷤ڛ+���x�LX|`$$�6d�Ϝ�f�~�"ǋ��O�kn��R`����:#[4z�՘��N"�*>�|�L̯�*@�|n�rŁ�쯨�*�z���c��$�Ђ�������%��u��#+��H�g8R��bN��-�с~:$�� �1t5`u�}&H��ɮ����q���7�P0�1���/�9li�A��k�T��|��e�n�^����[V�Q��!3�mqH0(�Myj���Ţ�z>��f��ۤ!��}�U�
3����j�kWK�c�+�0��1�V��u�W���Ls�)���'�8��P폿Z Ta��X�6��F�s!�y�BU�=�L���7��6^��[�A�] 7�G|��kS,VJ�ܐ|;${<�y���=ʷL���0E"UX1+�Ğ�p���7WK$�SuO	9jo�B��s '���ͱ�ɳu�T&"�Jʮ+�)71�Wy�|4�3����o$�5���U-�8.1�b�_G�+�@�|��n���AE-��1/lHhĶ�Uw챁B��(�	�pX ��RIz�wL\� I�`��!r�0�����r��w�@�N���" ̵8�JGǩ7�p�6�]R�	;.j�/i����+냀��-�I��t/�*�d�Wn`"�<Q�=��'�yu��BO�\��Ȥ��:*a6Y\��f����I;�&k1eòʴ�J�8 ��8M��NM�/�9��u�v���bظO��PW��c���x8�SKW�M�P���R�>,��I�C��9����ji����8f�R�:�'Pڰ9���	Ti�"�����暖(@w�d�٠��y�a���1عg��sK�� �w%hv���<�G�('�kfN�	#��n�z��r�	�0�K%�f>�9�
���"�&$u/�lr%������-B���h�m�iB���3�E8{ʏ*O���������q$h��I��, d�5�^��������L��)/lꌝ��Kџ��:� �s�l��'������O��a��s-�� y�(����)N^+�6��>xp���4�Sj�7:�0�=��ܰ���rg ;���G9����{g�&J_{����z+�� dC�w������,�y�_�=�o�39
�YJk�:#��Nxh�k��AS��n�9����~��0�ֵAx�K&�Aтb�H��\/���ú's@O59�2�^g�7T����J�Z��t��
:�Q���KI�:@t'�C~�~7�!��r� \9W��3�' ����\�n��C�h�FQ ��yy���v*�	�����t��]w�~_|��[e��gx�>(z����ߩH@����R���g�ywx=a�bY������<�fr&�' ���D1��� �%'i5ۭd�*��w:��m݊��	12���>�/��r��i�A��v�X�ꕢ1#d�G�-#B�>ԡ�u~V�V���0g4 2/��*���0�% �����ߓ}�3�RF�i|�ï���i�	�:��C3��0D-M�d�טG�}7����7��FY�\!�
��,�V�J��fk+��z�{��9�]��a���Q���o��g��K��m!�n�u��!& ��5*���͓,�>�gB�H'7 6��ݳ�c�QNf+�'xc�n[���씽�4kV��$���ԃ{��@Uǀ�5��c�m����=����à�;(M@�t�D=Kq�<��=f��5���N��?�U�tE�~[b�]����n��T�dk~�%n\;`Y�X�Z0�OL�B1ǫ��껥C۱����	�3�@f6�W���y9�emk'�2�\5�5���L�U�����C�fz�������i��&.t	S=�&��C`�����B���	ay����L�q�&V䞦�l��D���9A��.~��5iQH�9 �<<�~����ʜ����+pA4�q�W\��q����D\ۋY��4�X��^�41l
L�hm���>.��^�+e�T��������+�������͍�s�/����7�� �jߙ-t��뤅*[�Z�ש���-�c��W{�l�j\���ǈ}ut����4�8^��T�(C�9��o�Q��8�]n���g��͊v��S���	�lPI)w<��魊G)�`*��\שk:���K5���CT믣iT� �2��+++i�8it���k�m�xN�Ѷ�1'�p�S�,�K�i��)�V�lpo�Ke������[�R�J13�2T��圬��׳�X��y����!	՘}�Pv�PkI�&4��m������C�U9��\��(�{I)�p&�����w���� {�5A��~�� ���X���<��;�I����5�����s9?4� �i*�͉D���jNG"I<*>s���3iH������'�3�Gk`W�-�� I��w��bhf���2;3�tT1����8�D��4�':Q!�P�X���޼��b3�ރ�[��,Ƒ �)�s��ȏN�⌉�Ë���o���)��Z��5q�I \�Q�Өsܗ�"*Ú}�ۮ�HĮ�EM��ѝ�o� 2�uA�r�`���O!ܕM�Zh$��un{M`��
��6�iË�T� w��	�j� ���v$��Ie��?@�������v����.˘582�*т�Se_D*���ˌ��^Uvq�
�T��N;�g����k����	|�"�R�jO�/:��/Τ�ϯ�=��7��,?k�<j��⃁�z=y"z����ssqi��d$Bf�Jw��\�M�]ڛ�_a���ń�Z�ڮ���|08B,Z�$W?��=��w�g����rm$m��W49�!��� L�Ifa��,՝k�Aw�5 ȅ�q8�w6���o�0�؅��F��@
��8h,�5��(vq���j9G��v���R�e���[�[�C �����i&+~#��=�o` *ro���Х������5fR��e�#�緣i����wz���г\���|w_��$z۷���1�.����A/�XЫ�K�?��r�)d/N�>),v��^Su7J�]]
{�H��(�(�T��ZP���0$ӏD�}7��&������U�[��2��6+]ơ�>O!2am��kn�S�!�����4q�m�g�r	����
���9��рq�@��S�|�Oo���p$HJ�l'88l'c��̘<����&'pS���J�m�_�+�ѭ�ގ8Y��;Wb���덽)�9�2u��I��B���mO4��>0���q��-5 ����H/V�����!�
�����9��#-��c���7p�c�k�/sm�M�M&�s��7���������_��4\\"e�YtA�����? ;7������sJ� �Pȿ`��|V��3�������bx�˽l��B�"��g�O��Z0�j�H�>KbZ�q�qw��ꁻ���/�?�r���K��)5uJ���`�!*��}��?+g~ 3ȖUr�Wxɂ���!����n�8�_в�?A���&��MNS@��*�w ,�w��RX�?���t���C�`2=(�~֙������������?>ϰֳ�o�w�-��S �;hr�\S_�w�!ˏ <�Q#��o�ZE�/�`���7t��yO6)�_0�M �(
8K|v?^r釀;% L%7���?��1����Ïh��_����s������xBa�@���u�$�k�U���]����g�@ȥ} �K���n��h�}���	�Y!�S�����n��ߑ���� Hʿ3_�u��3
�������<��[ �֞�-&�Eq�� �`�ޒ ���)�:�ao�A���<E%o��ք����~��	��~11�ק�D�Q>��6��ۗ��E�J�I����h�GSKr} �w�A��)�K��ȿ����.LMMuʍ�C�"$o�E �}^�?m���x��@"��bUǢ���ǲg�~�=���(`:S)�������t��U`���7�3cV��G߿o���K�X�ŉ���ֈ���oA����	��T,.��Bp���r"��J��E��K ��:)���4��#�4#�O�yU*~�_\�r��Z���%j����6�4T�&�yo�(70�,lv�3�G�3����:yi���ѹ��N�8bk����s�.m���_ڴy��JG���Y�[�@Q{�'@�� �m�M�@�#8���3O���T��m���X�Q`j��'���	���r!��r��ե�v���TVVbc:C���N]
�S �0�e4��p\G� 鶎$*2��	���;����<B�}e'����O{#��ͨ��}�.��p�jM�D�P�	�z��^Y����C��)p8Klj���� ؿ`�ߴ��*�����j�S�ɔ�(�Iy������2M���PK   �F]Y	��#u } /   images/a63a4c90-64b6-4a83-b635-c920396f8e2c.png��S��C��`�S\��h�@��R(�^��w-š�Kqww+�B�������G�W��9�=;���>��9�������   G^� �\�� a��_ڊ�hV�ʒ @]<֣	�{39ue ��	 @�  �������� ��1  � �|�nS�� �T���֝t{���$�� �"�����&�/��M^Y����~1�<��IMϵ�'�	�T����tתΛ��;�6.+~����������$�at�� � 3��5r�E&N*�m^�'�g�B#��eZ������J���q�����i�r�k\�ۡ��*t���io+�Se�������֦ݤ�����'aJ������������F�!��T�5x������l>gP��m=�*�$eTɷ�d%�L!R(2��!�c#��т@j �M����������)C�h@~dHI�]��	F���>�/��C͓�Z�Z�@�x~-Vڦi�p�[�����?:p�Mt�b�t����=���x\�;��,6�������'�>�z�2�b�B�.�5L�nK�%�^F֦��h[��~bg����T��1�i �[5ӈ�ZKHUr��C� %��
�ѡ����ܓ������n��B�6��Pݏq�@Óx�y���ҥʢ�NU:"Tv4,Q1�T*�:˖�G���/L����ZoWB+)�M�00��&���-����-=$=̻�]
�z�XЧ��l9���Hp�f!S���BP����{�=��Z�ۦ�Ŵ��
����g-\���S��j��4r������x"���S�wnM�o  |�o�a�����x��t���Q�<��M9�A�7�-��i�4	K�W�DF9���o:$�XD� �ЁJ0F����V~`%-���'!���}�x�cp7!�C!�7A��0��]�<{�z�7H<<K�cH�'[����z8���%@p�X~׮y��9�NfL��N��$�B:�����|][&O]y�J�<��\���F�_��-3w����a�i�ʧ/��b�*���c��<Gh04����ɜ#@��u����R�W�
=jj��=P���B��_������2����E8����[Q������>G�S���0����~	Yg|p	+��tQ� D%)���$(�,�"����ۉ�VQ���
@O����`�C��Ќ�U��$Dr��f����UTR���(�V؁��9p���x~t��Oר&+댭�����\ @�Ё�F!��B�PȚ�[��pO�`��B������(�a��Ŗ���6��15���l��ꃶN'	���ރ}���@������q�8���\R��l��M�B��CND�/$h��E+��=��dHqcwwr|�������a�9�K�����ܻ� T<*�"��v��O��!Go @�\�-	T��Ң;#·�-YD�>c@��K�9lLu0hz��Ȣ��ݏt��(	l�m�>2Zgs�z������)�d�l��/B!d/+�H�Cұ�a �tK)a�P+�%n��K6���?��S�p��'?�]]�y|x��4���.w�b/��:���o8����登�~�oq1�8N�}ћSde̛P-y���LUF���U�">�@�RD�.�,�S�O�N��C�q"�t8J�;޼��0�-������kE��)H&b[JŠHs�	V�:G��b��a��P���^��9�;����9�-��y����9ص�>�����8�����w�a��lt��O����}�5�sKq!�2�4���i�Y;ѷju� � ���J�V
*�F ie?��P���t�~���g��<���ј@#b���N�T�.�@��V`�	A�*��&Dx@r�~+_\�>���3�� C�Q��ϊ�ɤ<�iq_vy���\������;��2]1H�kyA;׺Z��_��!K��, &z���R��m�3UD9ȉ^�����S�U��2>��`"E�]wK}ľR��k=�
�)�V�'���$2�5D�Ģ
�G�ƈ���77�̀@�!l�CX'�$�Z]TF��W׿^�M}o�â��c��� ty������=�V��y{�tvnO6TR��z�ܧ�Rl�W|�������	٪
(҉���d�"��	2u��޿�N�k�aY�Z	��ֺ?�O�_Q,=�/5wv6F��ߟ��&��@G,8ytdT kP���>[�s�^<���������=_�����6�g�+�U��C7d����Ʃ;v���#�����mI䅓��f\7�Hwe�|93�Z&�Sn5����U^렚�����C��Ղ��j���UC̳�B�����#��ɋ�/kgdK�RHL��$FJoF	��ATc�a��^��E!�1�d���W{����M�~g��iY��\/���^4GT�,O�[w�t��_�ϳc�.�_�wC��z�*����p��y��ϓZL���'���Mw������~B;���c)���Ve`qr�G0И*�}YG5��*����� �M4t�Y��b�n-�w/��SbX�2���u�~-����S���$ #�A�3�;�
�@oGi�a���κ{ٝB�g����O��Q��?�=�����}����|�8��~W�Kq���ز�/�"�˨ؗ�2���X�,Z�DNk���4�͊��K1>w����S�e �b�[+oդe���gLr��Ќs��\[r���Po���%%g�B�ȌA��,� S$�g���#(F�
pQ�' _����z�Wt�v��?cOM���Qaܷ�b����n�� 9���u��{ξ�4���^(|�-����&��w�OO1xY�x+/|���~R�&W�ʩ���<�`��<;a?F�|\��!��~�_�
�����o�����3�П���:��XA<G#W[������F�h�FI[p�0�ܾ$D�����r� 榘;���Puz���|����;�|�@���!�yevq{} ��P����eͽ�4�I~��E9�O�X�ޯ2�5L�$I<ؒ��Ff�$��
i��e��5$fkC���S����U,n���\���4�E��oU	�<��R ��r��[� \��X`!�S��Y��@$O�ki�"$�e�1��'Ԙ��!I�g����7�����YoG��s�A\�n�>�1N!;G�����CN�&�k�=���~���U��J��}�ueI�ohy���2%r�ks������p�x�s�)9Q�� �*����(�FV�Z�:?�\bn&9�Y��,4b��Ƃ@GA��ft��$,��sNq;���2�zxM�����#}������U�)�V�t�_mؽ�^�Ihu�^lx��떞v�:|  ��wݝ'����t԰�o�|>��'c�����=�Y�~M�K���:Y�q��Nw�+9R��_�}��R�p���CV�����=+1n㤭���]�6����9`\�o�^8�5X�n�vH�i<L�����	�'��EA@� �^��8�"G*�4�,�c΍�Up%���o\<�pN���cOO�un:c��<��q����C���n��ް�iOҭ�OW��'�q	����U��>�TQ�Ո\��BB��!{�i��-:���vwT�?��]8�|[WI�yIz��E7�'甧G�K��^�1Z܈��l�׸鎎4,�aHa�l�%)A�<��J���d���-LVV��^�������jg����ͬ���?3�|��Aق񝬮>���c*�����4c����kZ�B�a��!f� Qܽ-iЋM�F|�����쯊��Ow�5�y-�\�F:T�_�����h�%��_����/9"�pB�U)A�P�'_����ú|�������]H��b��i�Q��ꩳh�f��ou�M^�ƏF��E�.S)�P�>v2�)���B$P+H�d7R���l���P������ŝ�9AQ2 �I��i�j0�����(�T�Ϭ�ʅ����v&k7�m^���G��{��{����8(������&Dv����|e���W�|��_c{WyTL?����pL�U���2��}���Op	IF�@�A`ʳr�оvr��'q;&|I�.����6�
�,��n�0���N�>�oB��Q�B~�F��ÞV���HV�f�I��Q��>�zYf((� ^<w>����t��#/���'J�#b٫I�~�A\l���]��_�o�x"{:�z���}��1VYC�|���t��y@[�םo�Ecy��bˋ��t٪	\s=zp^kT�����
k��խ���Ev�H�w�i�w��a���?k��=��3I:D$}n)(���É�� �N�{� 镡_՞��k
�XGL1� zE4�`�Jӵ�8��Pdo�ǐ0 x��떩�Vy{Gȕ�����ÿ�i����4�X��a�$%VF�}��w�`i@��ʙ�3�(|�|]�B��Wć��:�M���z`R�g�Pd�.�>=kI:ꂣ
7��˷e�,�/���U�;�.`n#�N+�H�{�䗾6$���F+6?�آ�����P���}�to���.O��&��+�ɝ����G�ZN��"z� -#��jy��2}n1�f�G���q=�ۻ�h~����7H�)�,�$[���Mɵ���&����Fitԝ+��]_Y���3����	 �'����W�k�sT��c�L�9_��;�%9ΑV8w �L��>����F���΍-��+�������[@<��&����W���"xJ�Sk���*��E��x����Ō\��s񊎑aK#���aod���ԅ���k�eY�-�w| a*1݇�$�G/���������ԗ���g��g���}�
�t�}s��Έ����E(%���+�3�OV8���V�O���C=*���{�gȋ��eX*��ψ�U�Dc����M�hR���dE�R��o+Q�U:�W��Uo�/@�hfm3���-$d��p��[�hm�((�g��Q��{	G*ZTYL�$i��.U���}{��猢g�] ��|�_����#��ڋ��?t:�WN� '����/*o�k��a<秱��ͨS�H7w�y8Ś��v�&�H�tĵ�$�9��zS�~�Fv�݀2_�������'�d����n��K�X�����E��m+��>^%��RY�wq��؁f�D!=�Ry=J偘�4,��ʵk�Ʀ�U�����$F����ԧ	-I�u�"V�P�-<�Wi����<�^���̀������@\`10�M�T��V7 ���8F�ҧ&�B�$��C� �����A�hIU��/��E�ρ�;�D4��^��`�H�> ���V���^�79�\T�s�P��z��vJ��˱ܰ�6�G5�� ���ģŤq���Q��x��	rTC�7�g_��Ȃ�tF��\|�Y�",�GU�0tF�M+��^?C�t���B�W�$  ��-��e3�h&�I��o��@��6��iVJ"R"�,z,4�N��	4+[��g�3U<���Z�34�;�}�͔d���TOu��h�:̘ʁp�*���`�������kv �airs7,�̉N�9�_�/�o�'Uv��Ή�M��|ݟfYr��p�vz��y�M�K���`)�"P��MCr<XӠ�Ii��ѪJXyU�m���;&��J�qQ5��Z��[i7[��c)!�Po�}���O����UpKf A��0+�TU�I/B�C����j1+{,�һ%�WA֒�}�|����=PZh>eW2ݰ bH���@���M���!�wv�xd��5m�?9�xblf���W�cd�7 .���﯊�����y)�\{���(�t�����`T⬪f��(<�<����H�%���9�t��j��B$M�ilh?�ϱ��g��J,T��@�+�$�b�/���*���*���D���xB�eB�(��IOuChMH��K^�T��݆Uk�,�C!��%C�w�����{�)��*����.Bş��
���UUX!fb��F�9>���Z����j<���t(ș���h\$N*O����t�B�j��0��>~�%��O<?U�E���y�t�f���Znz�Su����y���b8�+����蛈�"������E���`���>ǝX~=���!H3�R�:���ќhb>�_eh��� &�P�Y���4Eyǽ�{��ip�>�(YPN�o��T��e�=�)����72,T&7�-�V�W_� �Z���ݣ���~}2EGf���[����<�w��2?_�y�t��|�|�����ί`��o�a�	qnP^��es�*w�fe=5���͛�� R2��BS�S�j��y�f�:��⧠�c��SئV��V�l�>P��_�l��Jb� ���cl/�D�>@*��+-g��v�S>�<�-B�2��S�qU���@0A &S۠�cB��S4�k�Y�GE�d�u�!7_��	.}:5��]�!�*�T�����5���Jȉ��\�A�<��[��m ڛDh��V�x��+���T3�f;y?a~2�Pʛ\j�%���I��Cb��.��w�J��F�c)sڸ��0�m2.C?�6�Z�S15�y�s�vp�S���v��_��]�Jl�����z���~JF��EE���\h@j�^!'��Ԩ���-X ���)0�aT4!-"��$U�U]���v�b���׷��nI���X�kd,���g�7n76��k/�j��hV�-e�`��F�%��UNĴ�����i�i�ՖB�& ډy�/����4�E�	����~�����N�f�I�%E6)Θy�N�j	s���ET�3��/EA����38� �LA��4�1�x5��`ʟ)��#�	X%�(�Q���i�}���Q�q�'n �o������gC��a�v�+fɑu�������O�Z��N�������Qc�ergt.M�)�K����n�q�q��e���Le��Z/�����lV���%��aV�Cҷg�DfU��,]+x��xұ,���E�����?�Jk��rk�������*����~Ù�d�q@�Zx�9.!�qʑ�� ���P(8Sj�R���{ċ>,U�G�W�~�j�,�a���ςhI_uҾ����Wͦ �CP�֟�5��o*h���{2����C��� �N��Y�z%L1jޏ$жM��qi-�d1Tt���C�7�8OM���Ϻ�Rې�?P�dQ��:�	�5��E:��O�we ��&)��Mk��?�4I(�i��S>���N�>u:���-lgTy�=>��>�_|Md�l;^�0sd�0��d�@xd�|"�U=$&B��["��v4���2��4�r��/G*)4	��0� 4�����(QDV�F.�fr��ڳ�H��U�؛*�%'�ؗ��}����.�$�P�i���q"(���?�&��eP�\����Q��l](�4`q��C~���O�C�~o�^��c�`�/U����N��"H��Gg������������+�tRE{8c�4i�B�0�?6?p��+��ַf�dv5�Tǰ�L����Ҵ�R<Y�]�7Ԋ��L����|=E,�����0U��:T���]̿l�jzi����}�"�y���d����/�?Z|��ix�����$�n�_ �2p�B`��kB���?������_���ud%�[�o9���9{j����OS���_)OG��c��2<@��/�`^t$P�~J�$G�#�LٗeEOi�2��D�Kؒhl���`1��S����0�v�!�e��7��@������u΃���ĳV�qS]�h�O:c��=<�UyT���5�P�����J�@�FE��A�F�5�'1�WMY��l�$��y�B@AuRM�<���i<��i����e~W�_����
T^��/�a���Еc���S����^���CX@���|Z�*��[N�MX	���?�8&��2�J��K��qX�����8��"���1*����]^�d�)�� ��}�v�!�:)����( 1�w�c�,_佡XG|���.n��B�F^��$(�Xo���ZB?��*��6 �gr��hwiC��T�LN�4���24�b�L@P#Hա�n�ca
�sPe�V����C�������Q�f�!עM���I���ٷ>
���m��-�e.����	2�e{ D]Ʌ�;I	��5/U[�χ�/>/�9�;��uN^[V��=���[�]�V;��OZ�ʇ�i���ģ�&R)�У,i[6�cߜ�
�o8�OS�1���p(?g�w.�V�x��5�VZQ8��P��Q���^�ԍ�&�3� �L��ȡ���߃5�?���%g3�҅F� t�u?+����<dݥ��J�<��YX3�x�5I[�bя����ϖ�~*aS��~ѡ�_� �V�a�8j:�v�s���5���!�ܧ�R�aGU�@@��y����A�G�.�鮲,�,$�H�Z�<�d�N:T��$h6������$��)�Fq��������J�C���՛� �x�g*�#B�Ox8M���3����@`ݤ^7Ni~�;�LeF,���v5$]aUA@{��y�u��`�0n@ur���">1tћ�ʛ_L��pP�[�)W��t�G����d���/�]�T��t(���?�5"��%.��:���Z�\Pi�K=�d�#�5��a�|X�P�T�=}FKɾ�s��w-�U��1�C�s��4�s�)x�5@T����O��m�g��eT�%��u����n�c���%��e9��jG���S�����'J|5�)j/	��3�7؂":�>�D�����筀��x���w�l�����l[���k�.S"�6�}��4�Ĭ�ek�d�T�}�v��.�.����ɶ�+��tɬ�V��U��j��A���w����T.�R�B�+�Ѕrl����_LE����(E��V�pև$Ʀ�_D�����j	����5��.=|���3�X(����զ�]C&�e�d֙R-JR"���X<v*{������c۬$��0�@;3�60�r$mYD�*#D���<R1��4Q�|����U���	��8��PM(�%h�}��B�?����6T�j�K�5������n�oh���ޖ[�L��p�W%�r������ �Jۍ�����1a�R@fv����'3_@��^���R���hc,s��g���N�í�S�n�4�O}�K,X�}x]m���*��q��X�'�$=��q���y��r}W~�l}�'�3�&�=����Z�GƎ����e����^$����2:c� ����ph��M�˧_�[�~'�[�Mۭ}k,���0���c�;2�>]�]�l�Z<.�m�<W�����c[տ��3n�~x��p����ڃ?�DL꓊V39�RL��&b�T(�% ��F_2'�E�oS��=O�0w?L?�u���r��u�_�'<�����팯�+�3���'�Y����s��<�TPt���������(�n���д�-o��Z�.Z|ҎdbC���u�>D���<BY�d���p$Br'�'�+o��_�K���/0u�	��
R'լo�@v���.z3��@^�C�w������ݝz�ʁ���-ˁhox?��g �m}��.��L��������'r�/��y=l�.���y�������ܦ}�Ik�1E�Ų,a�#�A�z��daL�Q�$���	��g����
��L0�<��7��_�.U�'7L�9��;���'�K�����L�u�6�7-���G�Mj��V}����a�?1E���g�q�:V	M�aY=}�J���.Z�	5I�u1HV0h�7ّ�7%�7S�}UY�!b⛒����K�2�TL�E����h�G�WX����g
,7�Q/E��@7�\>�>��kR:���s��M�42-�!��P����N7	��0Ƅ>�ʻdj��T��i������T�\����6��l|�@�w!8(P$��s�v�b{U[��-� ����MÎ#��*�O���h�97��]����|�b_e04��3K��hX(CYǋɳ�qQ�"��J��"x[\��]�*O�:/��*r��QHh���p��#���}m$|RWEia�`B*F�֒d���5�ɬ�����x���I��n2��UFw���آ{*ko�4����������^g{�5�S+iU��W(pH���R��a��'�,��5��y�����r�#�L>�8@�� �;h`�:9b�w�Y�kK�_����g����33�o�YM3l\rY��滤Bd��lGF�'�z�H�fhT����K��pX�B��dy�>��/
����N�����Ⅹ�kr��sW�h����w�Z�1�X�;)���h�jw޵�{�6'���0�c[��0���6R2��Y'�Z�w<��쪘(.0�}U��CI5�M�&�,z�Nc��x���ԇ��zDn�W)�G�l�.��5��b����ho���{��r$-6"v�аҝ�>��f�(��q{����H�y2�J�B�w���1��g��F���ɰ��X7���M�Q���QN�(eb�M�{}M������:��BE����A����Ȏ�1��9��p4�Ղ}��F��-�-F�f4,7�b>�'�+_k����4>kc��D����;�Iq��*�/nv�r�q�`zj�DW��76��*N@L�S���c����˩�}1W�����y����.ڸ�����\��ۚd�:���]Nlgƍ���r�� ��)z3�ҼIv���nӏ�� !D��˛�c8�Ц���hプ�y�����V��%hj���<L6lܤ�~Zw�g�Q��țp<�X��E�����2�HT�c��C,�?!�q��G�4 ��KPY`�87��C5C��/�_s��۾���V���t��g��T9�3���+�証,q���bT���D���t2Y3<�Z�B�S3!�N�4��U}��5����g�b�x�wg����3�ðB�}t1��B�,�W��ϤE��ג$�
A�ڪ~�����,_Fu���8o��FU
��1,�j˃ڵ�r!��D
�pzQuʭ( ��A.����*L�W�C�(�{�)ERj�ߦe�հ��ΐ����cn�r��J�j�I�:'e8>�L�O��x��fY�9����/�P`\��^��&����%�SHH�9�	:�T��Ua��	��ƹnU
��a���<��d�Y���3�_9�����v���i	����K'l���aZJ�8��ө�*��v��:+�8ٓB����j�7vY��H��l�+��Ho�1u3�����uUMԮJ����委_�v'�j&_��yt}d�*�~�E�kg�%�o���l���1��e9c��G���V9BD�eo�+C�79^���j[��a���1�|�+ώ�o��Y5[x�=Bx��-��(�����
�J�atp�n�yw�@���H���(+�m:���&��k�d��*[2h��$QX-*=\A�}���ԸtL}d���XY�URlݧ��5ˢ�,��K�}�.K]�����(`�����~����0Q�ң��է�	�xhd�?WD������YHf����Լ(�~++K��N�M5�-řy��C� +�u� mQ�x��"?���?�"*����T��@$(<�<��ȾK�;2i�q���P-ѼUJ:�Ѫ�!���� �k���hr!��b򪘋�;�*��ѵ3��9F�5��r.��M��]�w���0������V���w��5ڲK�K�Dq���/4_��P^I�NNR�����p�<I�j�C�/ʋU�^�2Qx۽{���J݆=wro?|���hU��#8s��h��er&���ƒ��1v�>�9��Ft���8fŃz(<�̥od�F4e.��O��F��Z@�I����s���҇�ύ�H�B��4��p�������ֳ���]�pp| ��mQ[9�뜝��=�G�-����$1?l��`M�b&I�<8�ÿ�uAׅ������|�;a���s⨵��ݖ�d�/M��a\7#E�E�4�U%+}��ExS������k���>���k��{�qyM��y-ю��4R�-�7�-�=�0n �'�hT�~�s��a�[�F��4Uަ�c�K8#���(��^�{KP�V����O3L�l;!g��i�� f����N�'G��	
���5�� JI�2�P�1���%[ �1E�Z�$~)���A������j9��o>���͔�M]	�n�O�)V99�
c�Ԫy�s�J���Aqh�(��MK!%z� �E�>]�� ���ޫ=��%Wr�|�AG�(`��4�᪈��m��s��)O�![�+�����i3�H����ӭL{���!��-۶�%.L2�Mh[��t���F��u1t�4A���3��=ߞ����;�^��W�	1��4�
*=<��.=�&ac1��L
=�l�eW���\��#����-��7t��ڑ��珆f��s����q�S�:�hE��W�8��|eS�t����oq��r����sC���CU��Ͷb�P%>�>�?G�Pt�	=�c���Ͽ��߻Qb\EЎ&$��f��O���L��4�Vdr����E�zcq�'��S�����A��9o=�\�}���"������*)̴�}���Z�uV�(��[�ը�Yj'X^S�h";Tɗ�4�k�Z-���6}z�*�?�����N,;����?B�ފ�Mې��K`�����<<���g��1�~s��1��n�#å!("�1��Ũ��V����Ұ�q��s�Ph>�ȰBD��a&ʰ������Ւ�rb��YqR���,j�?	\=�[{�D��=_�?�rS��l���˽V����|��b�U���b(�ྮԤgs�n��@��"�b8i��2�!�\Gμ~`Ty�Z���I�g�j���-���{�7p�i�D6:X>K��`hHgH��� Fg�_˹����9uj�VM&��T�g�� !���T�������H���b�}O>w�Ux����M�Q�?pCl������$�3�<L�k���f������5��Z�S���S���M'O ��|��A�B��[�TQ��IaGq�����菓4!�J����Y`Ty���n�����~��85~�N�O�R��_��i�S�t�2�92��
�}{|wይ�T�= H>��ɯ���H��%@i�K h�.kRc�\���� ��Xt�]��$+�N�}��ma����"��M�v@�[m��X7���`e"�li����}jG�l��_�N���X�]�٥ �z%�H}���^�
ө�׿�-ڀ�:����<�y�	Qi���r��O�5��Φ��u�j�����+��My�<h�[XVb���������lb3T��Y��zyp�n!㠅���8Rz�Z�S�N�~!��q����%p�ƛ�8�
���wgV�����T��Wմ Fv��U	Y3��ws1XX�Q_8R0�B7�<0.<���c;W	�3ͯ�wÓU�Z��s䤍�!���wfl۪l�B��0�6Q����AŖ���T��˵��|�/�S2�7am!���=}�t�1z#y��I��N���X����@W8%j�3�s��G���Y�����|%���F>����8T�?��Y<o�̉��4����]}����@�LP���.���>��٫۹��u\�
�zsy߭����'�T3�y�)G_^U���"���%4���메��%�9�C�$�ݱQ���-!��<�)�$��ٰ��+.^���7�O������`�ĸ��ȀK���k�Ο���]A��V�����0�l�h��d��5&&�I�cě2Ѫ&�z�-D�j������IE�v-y/^�r���k{?{�l��ן����MS�$�����m�_�Œ�3�XK�����:�����/���E��3ȩ��(�A7����,B��"i� yN�(8�:�O�i�˶��VhL�r�^�f� yX*
z?/�a;�Y��IrvnK,�T(���Mm�;���$ӓ
-�X9I��'4�%A���[���3HMEiڞǃ� �PLlS�W�h�$?�B̴���XHs�|��IlU�e\�I���J��IwF �da�D��:x͙�\F�v=��^�3G��XI��G#J;�/��C;��[��@�w��WA��Ƞ]�Ɏ���	܃Rf߳G\�߄�-�_�2�w1�k�d6�,�5c@MK���I�?����w�;���+f���z9��E�}��p��_���q��P�I���r�&(5(����cŞ+q-.d���^��'��E��4����ڰ���b��s�tbW�(f#����S8�':낷��#����B����N��>���\;�}�tW�k�|U=u��u�4�X^Þ\��>��a�����)�*_ɦ��c��N����9�
�^}�sxZ���x+���4�+��w�閣f�!�:��V<9�o*�p��U'��M<A8�y�fɉ>~>�$i|^[�1���|0�JQ����\�������8������ַ��$���C���|@�WyB~���U��Z�:K�,Oʋ�5P��(v�V���[K]�2Ӧ�P��UoE{��3�����%!�J#;�2�����(�P��4�p�u�㭥[��6p��{-�Ҋ���_zq��Uf�*���[:�^�=K*5^�&$�@��(S'�Q~j��,����AW�#9(���$�!&*Q�8�A�{���N5�꾗_H�} X��6K���?�^xmR	�'�����"iUqoH'CK��c��n����6�#U�е��q���q��sx�QJ���	�5A�NY�ס��S�_���?�5)�nfZ����V�l���IS�Gb��~} ת�m)\���7�\��X���jer���gk��G�^�b�� \r{%h,��� ����OO�}��b"�B�9��Q�RȬp�N���1� ǧ7i��37~�v�1QC�m�"L�Ģ���pL[���hq�r���SB�O�Cћw}d�[g�_r�̨�~�=��z,A̸��K���
zE)�1��L8�y�9"dt����ygߪ��R�����mH<�qR�QRC%�C%��	ۏ���[�t�.�)�&쏆U'c'�׼��,7P(�;��$2�]U$�\�+-&���u�ݝ2{��X�_�������XU��أ�� ���a��Q��;S�1xg�օ`9	b����A@Q�ݡ�+��2�P=�R�����z�e��KZ��&��X����Q�|�bv�1��MG=�E�J���,�ڙ��)�*9X�Gqۋ�w���p,���H���>���tV�)J���	�k[$���d���v���Yn��m��p毭�!g
���8�w����<�e�!�5�U�΍��M�Z�1l���@�`>�E��4��w�d�g&~���o�5�2���F���>�J��_q�{�l܈���Ɔ�<5ѱ��
����D~7�b!o VY� ;�>���*��uҍ������K�T�f�q��m}��I&��dHݺ����	Ӏ��8e
=Ξ���@�N��II�!K>��2f�TuU�Ss��Ru�Y�l˦C����m���ߠ�,�7s[�75t�6��ա��ӥʅ�����h�`mͅ��s&�^�>g�P�XQw<W���xJ*��,���yU0�E�-�OM`���"��ϐ�'*��âW�Z��-�\��HБLKR�V�Y���۴��?�I��X],��@��m%^�]��a���2V��p3�Ưk�a��zo�I�|e�PZ.P�H���ܵ����x��Ȉ(���
��'��;��7����L��)�S�c����ƶ�� b)I"�:�XC�
�-)�X{]}�n�������J3N{H��#�b@,
��T�yEf*�Oͼ��Z�(�d����C����'��I�2<[����A
�i�{��nH]�u���+Xt����6w/e�R���T��*,����R�S�N���m�Z|��w����c:@�Pݡ�����پ�p?HT+�������˽vǛ#�����"�zO$�do�(���Y�ъy�$!Үz�zQ�1�)^�hW��sLn�/m*e����B$��41Y��X'�J����,����CW�ðx��׉��#����sĔ��c�� �kb�T���G��(*�M�~��t���pE���9�ZԻ����8��Ohk"���?Y _w�8\	Z��8p���y=sݦ���ݟwz\9�xpx9b�r�һ�? )@ֿ�+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs���� @�|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF� @�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+ @�Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�Ss%�-N4�&�ĶmMl�ر�cs��N&6&��[;�y��n�_8�V����XU}�ս�Ew�%_CX�d���
��#|hwmA���-$Q���g��aQ�!Vb�P�+��|�l���5��[��Z� L��V�ߊ:8&�&�� ����2�ꀵu�
ӫ��	�T��Y&��d�Z����rx�Z��c���㢠�;�f!y���v�����r��Π9��^q�ˈuT=/�wE�t�)�e���.���W6��{�pN��Ħ�`چ��S�Eq������6�Rט� �w��;5�����2�]�	ɒb<2__��J6a��.~�S�T��#�:(�`�G�{���&8�J�y���gi8�z+�d>�)�ـ���*m��k�{���kJ^d&�hf_��߀�(���q�:�B��_���3(��hx�c���Ϻd"�Y���2�!���آ3�H����������u��P66��ؒ�ٛ�$p�[�|]p����m �.�����)�m�I�l�4yµԣހM�����o��8.�0�T��Qa���X\�#���R�yB��w�瓕#�uz�(��<Z�K�v�4�wZ~���pȄy��u���H���>!e�{��3s��r|`��R����˿�����&��JuJ
ļ�g}m"�fP��������"���nRR��@�ڭ"bhm���3��������d z��� �}��$m�5��h\Hg�6Al���z�C���۪ �,IA�O.��t8�9--��ي��v�����:�CT�M����[��|���w�� !L>k=hx}#�y�����D�������+SN��w3��0?�߇T���I��b����ݮ"Lg��ne?̗��Q�N�����F��ǫ��įІ T�������A��@�с=���4YԌ'[������������}�gY����v��u���ῂ�Q�mр���=J?�Cl��4[�������I�B���}��p��8ݹ�����e�fA��"����,N��L�+ �0b��M�����F���:y�i빆�H�8��l��zН��c��!�0>[Y6e�肛P C����+g�窽�'<Ɛol�A{5ޔ����� oΉ�x!���]��+>!�s�3#k8*ꯃ�Z3Dl���1/�( ��TQ���O
�wk���]ˆ��ݶ�?���}s�1�j�x��Aѱ��|���� XGŵ��̴"^.� ��Z\�F �!8	��{D��(ҧ�Q�2�%D��fG��<D�NPpH�h�;F���u�yl_9?������G��u���c������g�tV�㤿�i������,-6����.�o���p�����%(��]�& �)X�\z��Lc����%�JZ Qቮ��8��8s�8��H`N��Vi1���¾�&ȕ�&���&�!�=�Z�S�,ĎJ:tKٌ����0��7�F����1��&�mo���V(��Ɉ�v�n����N�]~6��Lt�5o^NUU��!�8��c��.�����(+��/��9bK�p:���N\�ZSn���:� ����S��+�	�UW�o���"G-��Ѕf'�
�w����-_
`�7/��6�pʎ��>�Iϧ՗TeԥFF�"TY^/��o��j�olr��cWb�ݢ���\���7�%N.��ɫ�փ���;R���(�z<�_By�x�D+0!A�.}�$4����*z"�OU��¯+�_�GQ[��нO��YQ�KA(3;o7a�i/��w�ʀ�J.�`8 �S"v=KgÓr��T(E���)/<R�Ղ>:9`�ʬ���3|YRY�Y�������^'����{���9"��|u�B�Y�Z�e�����|�3��c�^�^P�����E��!�s��V��K�	!������'�>$e_�?���{�:�?(�=�l6(����h�&�|���Z�Ă��9��W�ֲ�I�����޷�M^B�c��NK���t��C�#�U���|R�D�{��eS��*���N�%S�m����Z^��X�v��<গ���1~�cKo'�����ңP��*���-��Y����FhII��u�~mC�/��S'k7P��R�U�v'�4�_ѹ��u�Vp��K�^g�)��\�zd[�Э�j�N����������
��O��J���-T��b�/Z":Mƪ�O
��rZz�h`��b5�r�o���jӱT�5�B�R̥a^!���6����g��2?0�_%	_1{p�9]�o#�ȯU�N�NkMѹ���Q?_m�U͉2��ʢ�~љ�8e`�h�rx�_��_�[���>g=?E���n?����}�_~r�'��|�+��I��K�4�BY�ur�cg�d�@�
f,���$9^�A�u���1ؾ-���i�M������tZ�활f���q���Z�z�����W\�qZ,(�F��N%�QbƑLiv�usU��v򒯡x��U�("`���y�"�I���%�:���9ۀ��/v�#���+���l����
�
�X.z����YƵ�C)pr-=�gKe/�Б�!�d ��B)"�� r���yz~B��b�a1�n,�"	� �t�C��E���e�n��/b�g5��g7�诵��g�'�����z��K9n9��m�<�`�W���5� Z�*�Nt�yXkz���O�5q֠Щ�X�o,��%�>W�uV�ޘ��/յW�{"dnA���s>DA������C�]Ϛ�S�+�+Fv���������\���T�?��=w����<"�E����J	u��(���k�g�ե(5��Q@����x�o>vN	��@�����5�n��#+�{�"❮K9p���5�G}wUm�L����l�/0^���4��kvސ��2�e���b��+	O���y�l_��CH�o�]k^jD'�i�M��_����¯��]��	��r�����j�B�_Xr�~M ���ޅ��<l[ �b7D��z��b��,��QK3�u��������}�`��X��Ya��VC�u��Vu��;�W-�2�k��1:����M烡��!�q:(\���T���(v��x_���r{k ��Ͽ"�'����g'|!\&G��\a^z��$�'m��Gߦ��3�+�RS�O��K-������ULؗ�"L4�����)���d�N�=~��˭ �P�L�������\��F���M�Q��uW��ƭ�5N��^6�ӏ,������IL�,X�3(���)�I�W��(��f��+=��Y�"���lAW��P�xߧ=��/��p#�������A�7G��-z�F��U�"�̶�~�K��^-#yD�fk���Fח��K�r$�\��:��G('q��k��B�����ڪ�>�ٯiL��z��*���4.���\��}/`5V�H�%��묇+U(}�A����m�w�7�3����!�g���M���3��&�4�,�^2B�&�Gi�<�����J93P=P H5�E���V2@?R��'�~S���^ :�ڄ��&��.�{��C���}�F�	���΀'��`��l��|���%-J����,���t7��b�@X�E|��D��ą�9p~Z��o/�W)�؊Pδ�)}�R-�cG���z�f�O� #o�����U6Z%�Ѹ�2=8�T�[��L;��t�8�pi>��X�*���F�Zo���?���q�q�Z~����C\�WP��Q9�T5�&f;jw����w˱i�3Wh�r	ж�����(�rq�NW�")�4�f����k\���B#�`���,'B�1a�M�-5�\lw/�m��t[u�-e�^��:@�}E^T�qo���i~m_��\?�Uh%��%�llfu��O���\ղ�h���!�\��L���ǨW�_�����x9mp��?�I\��|4X�]�����������,3�ù�=w��P�� �h��*ȕb+���0�����Pk�Q�q��4DNI-߉�Kɿc|�G�(�8Z�A����m �˷�8q��3D���`��f�~����Z�d]#hxi�G�թ�'�p�e�7��q��֚�F.��C��ȷ��+����e`��ⷕ쨲y���YP�-���	w�~׍=�,�������X��Ȍ_���y����F쿇ٶ�5\���q���Q���p�ǚ�*���Լ\o(Zۓ�h�"�n"}W>M��]M�^m��n�0��5-��{�r8�Wj�IO�י��P���V�H��Q?��i$Q�.ѕ���Ώ)����RXj�KM�P��A݄��D���G7�C.�(���F����L�뺔�l���ok)��]����EV�Z���L���|*��
Og�k�S�������jC��ޤ^�W"�$�������m0����Ӓ���@����A�⩍[���cr��On��E��K�G�G�E���[⚬���{{����ޙdM(��q�gK�W�F[�u-�%�2帘��L�ӫi�\=.�i������w��aNa���.�H���G\��9�3����>��a��M.��9�@v(e=O�(����1:uDN��5�B�͉ځ�*eNw�vG^��Į|(�y��C�j�V���U�v����
�l/�)߆LO��M�@0�����ISe��v�tY?+���V�j=x%�0%�e�oJ�S�*�!q�ƾ"ID�kw[u�t�ܵ�ڃJ)�f�Ŀ6,�|`��z���؞L��>|h��~X�\f�0�@��Qo(%`�����/��ү���r��������z�b׮�4��L���u^7�;ٟ,)�[ݥ�K��
���G��P͙�I>�S�5��(�C��h��OJ��<F�88�c:(��ܮy;{�c1�8Pϐ�z�2�"�䷗6&G�����1,�73g�0�X�J4�z9<ܷ`�����/�2
BI�Ђ��t4A�E�����gїw��W�|�*WZ��ز�Xax��*�KeI��!#�q�Xو֐����R�W�)�ޡ��+G�*z��A���bLC>�i�޹����Sa�5E�@���ƀ�Meٿ��9H���lh�]P]��Y�ۆ;5��-���)��+�P��=LIz�Cm@wՍ\�H�Ţ8�Z��'%z�_4���T��(�sU�R�mO�(�K��{��/����S�B=º9#nB]2u�$&D���@��&�U�ܷE��?)��y�ȉ�g�v����l���� 3.�.�r�sr��d��'=@�mi��n�	,�F�w���8W��*
���jf\�,�dvȂD{|�~\ �:�n"J�?���G�1_�ʆ�9(y�Io���Ȓ��d������I׾��%�@�J��:��P=o�GRj�r劘_��2�VBv�I<,js�7|�v�P�NU�����
(n�*Z?PG��
�����p������u�Z�H�m�� ��p��N��A���|q��:r��	6��"y)E�xM���`Ġ�,&.��{b����&\��QS�3�3j�x��g�Q�;��8T���z��~���/�\�������(�5��1���0�"����H|����,�]�k�aR��L��l&'�G� �c7/iE���4u����F��y�\��j��d���"�z 9�K��-�d,�Duq�ݏ�T���US�h-FiŮ&S��G3�H2�F' �^�HDT���ewz��`�D3�=����$^�i�9�����3RhT5��#��Y���`�+�s��ok�a�d��?�XM���tY�A�ȷ^9K�O�~��<qe�~�)J����	���F���?�v(fzT~��)��&�&��#���k�����P��z�=�´b��55��U���T�G�^X��6����[�B�I,�И�:Z��y�/�"R\/>��p�ai-V}l���8)��ӻSlB��&Q�~B�:J%o`���2^/(ͦ�dHМ��Qmp�����s0У�S�4�����1� ��+]�s���|�y�	�3�R���V��n�q�/f���=�h�j;�_Y�0K}\(ޗL-��&�m��~u7�����J������ȉ�[r��k��'o$Z �S�gf�Dˠ��B�����|yB۩�]�R_��=�+��(h�?��ğ,�7_{�׆�g�y��u��x�������MP�KK��h��K��"�
���������}�k�m|���M�k�
��s�Џ>��-�خ�cHH/G^��J	{���`ɠ��޲�8Z�E��YÜ]��"l�b��O��$�u�������v@�E{�����������jNĒ��\p����彘��ڡt��#l�d��G������B�ZJh4�������co+Q/'*K�T�_8�h.�#k'���`�jK�$^�}���U`�|I��^�;���=^��	����!g���� �u��1�Fe޿E͆�J}�0�:[�y1s���>�xa�[uY0�C4R��v}qs�R��g�}�;8^�W�p 7�շSN�z{���.	�"����#[�L(�U�R�*GV�z��ݻ�8����+_�}~T��(t��F}ެY��HՀS{ũ��6e\��?\!�p"%�[�FiAeaj�*�WE� ���qx��:��Ċ��HƮ�Q���a��@+,H�}�bRc`Wj�H�hH����l6��a�2!/^�Thc��6��O�'�����{��-�c�B.��l��:uk��� ��oGb��uL`�M�oW{ᗋd���S�2��#T���IQ��8�I��H�p��/�,s^���{��۸@���ɝ�R�շ�=�F-h\�#H�7l����&:Ky�7��2������:��^��i�x�����}E�������l	�����D����y-o�x����!/#8"��HL1z]�Qf[?E�X✙P�l9!'��`c��LvZDT1�%�c�$���2�i�Yٞ ����;p���Cu���D�QV����&?47X�"����%�����f� =Hcx��%�)�k<��d�:p����+Bj��Ƣ`������Z�;�	��E�V#�Ո�e\���"��v_)D��=�?qE��E]��qB^JN2���w�U�Xy�|��ț�����E=�n>���{ѣ"���������I5U��_���:.��HF16��w�E������ğ,�>�򘚬�
TtIr1:��M'�̛E�����~&�F���so��{m"��#�C��-��WAKt�h�ǐ�e��Ņ�Q�dRE�N���A	�L6�9]y��+bT&�|O�
e�>Ghi?Y_h��'F�R�mCInR�<B4A݇�Tx�]��?Y3�A�4X��J.�!i�4(�&�:�r�+��M"�(�#�1��{�43_
���9y�̚��f��8�2Z��8�����%>g@����F�J�E(A�\�­c�w���Y�b��$�G���(_SJ���N��9-�����-U�[ޏvI�t�6J���M$BN��p|��v���J6uM�lBH],5��N�w���!a&�r�����D ��I��Xm�2?~�J�t������K�$g}�;�UpG-��jN�'�Z�UK\�v���4:�)��$�JK?�8f���5Ù�c�3 ���vBJ�#��%�,Xjy65Ѻ�q�\@\�G�{�|��md������=�]����v�Y�����O%m����W���¾��Ҟ��My	V��![{���M���<kr�h�Scڑ�k�+S��C��<Q/�kA���Ъ�+������1��YF-�XUD��.\�� ��#�63���GH˂�5E��S�3��t��ֱZ�3�&3B@�ݠ���wN��$�v� C�����h�(�����:ל[��l��y�6SiN����M�3����co&U[���y�E1DA�p]�[۲��V�����nͿ+�x�u�\���H�ljH�}f����#���ӥ������rT��hu��j�B����=)N�R�����$��C��sN�/�&˳���d�~�e�aV����Jz%%���t����[�p!u�ʒΧ�-oPh1�C5q`�B�r���wi�vT!Y-f޷�R�ua��ȶ:0��5\�M����ω�
0��t����AxI6w3Ё�Q��ێ�������S�i��]���%��9��l�,���is$,�m;�m$}T\��D*�\���'�� �Qr��c�"�6��͔)�r����G�1M��yi�Y�~(����b�����+a�2xb������P���1x������0bw�c�ں��sjg3%���ig=��c�J�M���K++̦lDBHC�����:�B���1���%�ȲB�T�z�F����W�$Ԯ�.���Ǒ��i�T�&B�",�x���p!/�h�5r%`1���x c�{�v�)A�����u���j��W>��]��':�����Q'�eP	~�.p�7��^�p\r�K�HUAK% nzT��`�>�Z�7��'1�o�[p�s����/0��r�~����r�J17L�MTE�=�<4���s'�'�pea����$[��UA��`�"/p��IVk�,�̀��3 �ճ�~ %���8/iA�|���[!��j��8�w:�'[�E_�S	�`��!�W�Z��(w<��`;W��]� �w��ȥm�*;~����<k�l����4�}��%��]��v.�6�E�7�/�7A��G/�D#�ؼ�������:��~;:*�r�z��5- ���#f�z�t:�O/�<�]�����ӝ��l�"�qŜy��ŃQ�F�(�����s?��P���j�?F��{7Rjy��%����.\�jf�M�>���I�&%� ��Χ��׉I҈�����6�@�xG���57��U�z��nD������yu����+Sn��޷�[jJ�.m]^2�o��/��N#�D���De�(ʲy�2MY�E&����3l�c\���פC7�ҁ7��9�GH(�Y�:6��њ�ly9�vm����rFg�Z�|�OfP��f����t4G��n1�t�yݼ�y���Y�IGGO��{⋶M�n.ۥ�·��������FòU����C~���c������bI!cpl�oA9���(�P�68���i�~���ds��I��3[M-?��b��6Ɏ�\6�|�$���*ߖ6�"�E�����+	��c�幃 �wI$ 7'7� e��.�?6F�8�j=�&��,�yq�Vq�®!�l�W��ݠ^���N��gz��S�8��k|��D�CZ�R��. �
����q<�.[Jg�6�����9 m4�2��A�'�)����<�҅!I�x����>�~�!N�����g�^�>��kH�>�"�/6�X��F�:��iv9A�h�M�����u8��3�q��B�$��7H��/g�2��+�
Ui���h��c����d$�JI-cF��R�Γ��
nz�Q�q�n����P�8��=|���c����SC�Z�z�8��<�i�"B�����Xv��v}u��~w�^������LfK���OM�73�ϹI�;F�Ĕ�Iָ�C=e;BFQ�@�i�.2Q��ə25���:j=��=�r��Du�ʋ���`U�D=�y:�� )ѷ3y��q#�s�x�z���������ꭻԠ����\��ոHOcR�)��Y'���22��gZ!���ZI���쎓��ж����޽j�~y�����ڻz%��s[au��v�!�w�D�0TR�+�T���&��Q�����W�hǙ���'���݌������y�OV�e��W��)iϥ=�M���w{���CB�l#��Sa�u��)�N������2j�t���]q|�v*���RU�Tm,��AU[��C7	Aàu(���ߥ�೧���;U���K�x�?n�D�Y��v]	����ď�P\��C���WP ��j��.1gp�����&��)S�2�؁)����
2`_@�F�>ܫ��g��^�aC_v�����OJ�[���;�����?�d��	�����i�w��3��Lu���/&�Hw���bY���8(U���H/�3T�;�k��td(zEzӸW�tY^<���ZiQOt�Ұ�T����0������w~�њl��X(�Ob5m�jk�%�\q�A���y|�*�&�&ۓG��Y����)�3��fqH�m("�/�xӛK�x�{�`�Q���nƋ�������{Q���?����%�%:�r����.����HU�G�g�K��O��f�/&�OT���n��V��Z�+C�� �B\�VF%��������X
����]��>�E�Ӯ���h��9�J]h˒Y%�cݿ�S+h�3���8J1��<�k��0��	ۘ:����*�9�)��Ier-�r�xV�S��'���U�(�ʠsnwp�r�p�\�(_8�y��6�6��A�=I��=]'fr�<�RN
f{LS��`v�_><�@��)��\���Yx�d>JK&�����\��yy/-�l�?��V\�n*ȱ42�9�9����?��x��y���ԙ��H�q+�E�p�̓�+���q�l�|m��[l���������@��F�Tt�kǷN[MIQH\�f���
�G�v�~�wA̐S�����u��]�|����ZU
�s��ߧ�p��ǖ"�t���z���O���'���n���3	%O��2u��at��슗3<�?��U_���>E��C̟�l'UFp��jD�=?Zm>L �z9��T��&�A�{Ъ�C�NWY���O�3�^Lc?�	�76�f0�z�	�{�й2��C�#���#��Z5��H�	.���mB��j��CD�8?���鸔%��vo�� ������$�΁���m���.?-�m'ۯ��ӽc�gLon?���T��}�n����2B7OH�����;��[�i��a���R�Yu[~h	m���T>H��+}��Xr6R~G��-������ /����K�bǧ=�g�v*f��d̺�äx���^k�еW�y�JȦ&���t]��$�*�gSvmk�/,aD��W�Zۢ/�ϟ�k�7��+���'32����{��=V�b��/����?��/bj\���mH�U%����q�A)��=�a�����C9�{<{�5Iap������8�^��CI�NO�7[�^�����T����[dOZ��n@���gڊ;�J��bߢ�>a�����4�GV���7�J�sW��&:G�u�2�՗ ���mp�&nK��u�#�~�B��s�629�DsVW	���1���⋬QK���K�[yO�V[-���8mIF����E?M	�|g��))�P����h�B�^Z�jJwذ�ȁ�,B��9/=�o�N���*�s�;�!�}o��5_f���F�q���t��k��������k ����������%���.�y
L9�\y�*��+w~�]w˶���T�V����0V��.�33�H-�T `g�Z�u�*�n=jY�E@��#��M_��M=�KN)V��`~Ռ|R��wXN�3�u�$�'����eG��w=�@B�6������#(��,cЖ��N�^K��'�V�pᎧ`��/��5���f�V.��ws���p5a�"����~��b��Xy�iY�%�n��o��  �tIR�����v?IU.s�cmVE����X6�Ԙt ��ՎM�Ȯ��ݡ�c�,��0�-���Il��}��e2�⵬UU������)q͹��Y].�5�����?O;=�^���~Gf���N��f�o�[�m��8���NOW[ܯ\�D!vR��$!5E��s��^NS�^����	��'q�4d��T �Se�N]���H2&P\��쳔׎'�@܋�"���-^j�H�m�_B�� SN�9��Uq��DxՀ-���S��mg�*��/ozUI���t�V{s����±K�'����!���8��5l*3��<�Ep��2Z��}�8���v'z�?C���g_f%�N.*�^l-\�$��X"gÒ���І)�c��j�9��T��P}h_#�u��@��7�)FFMì=�N��<�T0ӏ-.�>K���p�� �lʭ��$�/����q�p{{���Z1��[Zp<���yˀ���Z�7b�;���ۄ�W��Y	b�p���Gh��?pBϱ�D�KJР۽��E�bضt<��oo�X�΃m������[����Qco��ɉ^@UJ��h��C^BP�QI�N��]�.L���LΆW��L�HC�9�D�?z��<�Õ�`�V�0Y�17�fD�X�1�k��\ |x{� ����ΰ��k���<v�� >��iF�!�ol�S��\i�:GR�ǬYֳ�#Ru��W$�<���Q��-�ӣ�A3A-́���\[��|hϻ�03r��@L����&<d��c@^���IW��&������b�V
*(/�~x�d���D���+7�gUc��խѢT���j{���:y����3o?�Zwg�[���p�H���>�_/��}�&��!\�z���O_���x��e��4�װ����|��k'�1\����h2.��pSm|���6�ɚ~�<$v .r�7_'�o�0:�nP�Қl:���1��()��w��f[R
�� >e,�e/�E=7&�8뜕e��w�j5��1�HW͕�Ӏq�<u͵^��Xz�c�}�����D�\i�`��!�3(�j����S��QU�z�"�E?>�t�<e��� (��Cak�#NK+��ud�k���ƚoIөg/���x�M�$<󋄧//����ad�!Ϥ+e��o��.Ռ�]�;�M�hz���Z��^P�:�
x��za�"v���{�]A�o^��Ȫc��6�l�)�6���ܖ9=u��(�:�Mu�ښ�B�����J�od���7Un�-;�$#�l�[C%��x��󲲲�����[&�Dә�-��p�L���Z:Ҧ�eEY�ha,gU�V1;B�G,�d'�x��[)>�?k�(f�2䭬�>��M��](v���|��-�Q� v�\�x
�뼯���U���/��������E��T���x�A�&��fn�f�g�b�_�`ca�ed�adeUga�c��c�ga�ca92o����� K������ƥ������������k�G���T��3�?PK   �F]Yԯ�|�] n� /   images/a794cf5c-4b1a-47ff-be53-d48f5d14bb41.pngLZP\K��%������%�����k��!����`�w_�����SEQ�5wf�����s7\YQ
��+iqU�%�W�(H�o�-$���\De�Q������(��C�����J]�%������������'www6+{Sc�Ol�ǂ�00T02��=2�==�>-�>�׍�՞��xg2��,�U<�W�"@���^����5!�%�;�nr��<넨�n��~�]z���!��ݓ
$r�W����R��Fޥ�X�C���
6}��t=!d�4�@r�7�-#���!������>ta0��ü[��'8Xi]yr��k�­�ތ�����L����c|�����ӟ�t������� <��!������J�}_�{��=�����Ds�c�����_ü��,5���kL"c��m������#o��mU��σgR$�� ,��f�h���a_a���;�х�2!�b��p<��jl���.E;�����ti���j9�_�]�'^1+Æ��ȪK��m%M��#��1��b����*���H�RL�=YөWz�\�\
T�n���� ���nǞ�����K��Z9�	T˛���2qXWŃ���p�e�T�f.5*�h��=�cPA��Ҿo�N�B�"A3�L�5�߈���R���Fq��a���4�"�1R�#c�,�����W֯�ԑ�� ��Z�꾝
Ne�7�g� ��3����Pf�3��Q%���a]�_b5(7��1���J�č`�^#���\1�|�d�^��Ex>h ���b0���G� �,=u%�
���/���q��-{�jt�l��G���S��X�f�L�'�>���Њȧ���$2!�~=[�)��ߓ%���/$6����]D���a@�U�b�1"�ŽLQ�j���#Q���х�6q)�o����&w�O���#�n�qT;*��R�����6x��0�Θ���b���J?E�d�m�Z����������]C���t���􁛢��wd���� ����ߑ<�b��J|a�RV��9u�6n��������N��tw7�^3���.��H ��_R�
b�>r'	�35h71�����]}C퀸�
�g&�'T�`|�_��9�6J�1b5�=B$��ƥ?�q7����ō5�Z�Ѯ�: ��ƬƱ�� ��m@�,���}�f1T#!�݈7zԄ*$T�� �˂��]R�H�T�e�D��B�	�G��'�^Ef����4�p��`N�����d��+p�{�t����L�ol�9.tqU�f�'�8>%���Dp��u�%]��B�0��ؽ�<E�D������M~��W��v�����L�����?PK�V�<�b]햫������Y���,^"��a���J���,��+�5V]|U@�3 �=?��M��#\��ʿ�VcJ��m�}*�x1^��O�V��Dܭ���y]���2m~�FՏ����f�8GԨK�Ƭ�eM.
ZxH�4L�a�
���t����G'�r)�οTl�U�l�/:ט��J��N`^Ŋ�q�f�$F�_X�$PX�h��n�W���ư��0��ߍ�F���?̰�5ʩ=}v[y|D�������r��oa�j/Q�Ɋt_X�mݦ���+?����x^�f��Rl���`u CZ�cl���n�{C*���8.�U���h�זP�@�2���?�2�Xg�/&4��9����Z��P��B9��˭���� <F�,~��Ұ�a`]BVݎH�;��cR��;oϔ<I���;�FY�:���!�{���Z����UF�C�:��n`*�癮��e�0\���Ԑ��\ �97��g�6�V����vs-CV�G����1W�i�)���ݶ��ܤ"���������onޖ2���p~
e ��S��������΄���X�D�p�+d�Bc���(Gc��B�b#��+��Z���F��a��T�ɡa�a~a�nʩ����͡��z�/l?d7t�4x�4t7�`D�7�^26���l*j3Lu�k*�]����43N�g<���In�|�^����=�	��.2��^½/"��\����&Gl����ܸi$wʿ!d�V|�6؈WB�a?��<����z�]�TfÎ���D��� `����a��7�!^V�e�C�_����'�`H��1�P(.)� ��T�=h��E���Vl���P���	 ���T�t�7�Tg��>G���P��ӉW!̸ �V�u�Pny%�� �w���µ�C!i��>������UV��󡟥��c�U�������J=���:��uԅ	B��ΰ��&���A�g>DŌ��:�.?�0;e@�\���Qd���d$d>b�.�39_��mqe�8n��"�n��?�?�檿�d�c�ۭ�)t�~���M�*_~���w©�{��M��pq]79��b8̕I���<d�; �ĚY}��M���֍qگ��4�r�R�о���-	}3�_j�GTP���^/��`��51wЯ��D��<��M�����hc�e&���2d	+�3j#C���!hS||����$I5T[�R�)����(���Q��."���|�B`W��;��1�z�dτ��c�|��{Z��2�CȞ˵թ��X����>���"uS��}'�4|(�ٿ?F�1|U���Qe5!�W��o:-�4[^�/��M�]����'O��\l:tR�cD_���"�X��I�@ޓM�a/��QX�"������m��f�;:�uz�3�b&��mEs����L��Q��6�~���Z��u����NЁ�qY�lU }ҷ�U�3Zhr�MP���~cK��L\ݐ���,��K�U�<�H�vM�t11�?9a
�]=�[�T�W#&u �i3�	���5[��U�dPPj급�?�B�/��T7��3EA��F�~�K�S&�S�<q�~��f԰U���[�bF���k�C����k�[>�пI�0nwS&O԰]oS�[S�L�j2�Ě� tޡ�p��Z)QRWVq���!0#:g��f8Tujʈv	�M͝�~�;[���C���/���f�ɷ�;��������K�!��
JC��(a���,hk��e��@'5�DK�LƲ��Q}&)�9�e��/����oOU����0�r-���=Rй�{3���lp��_D��a1�5��5��P~�a��j��[�,*����K(��u�i��
�>\f�X]IA�v/b_t���g=d�k3��܇�ý�	!s��
���������5|�T]m��������i�$�_c@��6�@D��R`���X"s1��X���HzL�gES�����3�7������I���g���WV�'�����&�	T3�6;ղ7S;Sf.j����3��U�T�/j$�Ai�]�1T�ru��6�ʹ��7�|��q��������ͩ_1F��枉�����](9�E�K��-遹e��*����8��.F����!�g�Cz
5q��0�mԥd4ͩ9ګI�����$�7�ep���z�F�EuY��_��i|��>H��\oI��ݚ�Ҋ�J���QОu���e�����%�/��"����zk�gT��/�w��1�Q�}�*�C����9��0��?h��-/7�:�0�~�9��m�,�W��%�"�)�I(7��2��%@/�;ʹD��m�8�j��C����M�|��`_"�u�#�����9A�-H�Ẃ�x�)L����8Q��5%(e��_��4�3ſ_�ͤ���>*�n��7X�v�����eN����nQ9����yc��u������}_�~����P�D�p��i%�Rm\V���F��.�K�c�h��ٟRB7d��\J)!a_aJ��,�&����9�}d^]\���0J���y�5r���b�|si�@�_���6,�_�T��?~��U�0����!���%Н���ԝaR�i�+r�1ڏܼ�����,��T݄�=BћOצt���!b�ʫY�@YUl��i��c�,Z�/��;�/�p��Y���^�Q}ZR]1)1����cG���/:s|.ӱ�޿b�����Zo����X�.(3�1�$�m�d�߄�?��yf�Kc@�,�����#�._�e�p����]�~�E���/qT�����n��ps�z���O|ۛ;�Oԅ�H��Oꠘ�d}��rh*�8���f)�U��Gjs^z^.#@�&��[�^�/՝�ɣ�r�}�Z[`������$^��3N�I�]��2&��3��K�.J�5�󒔅0}��lSŒQp���.E�� �l���#�4fYh9g���Y�����{��o�wz��z<����eHaA3�kn�_Q����g����oV��"e���>��HjK|/�r��rv�a��z����[��5�R=o�R���:�8v��i���g�(N��!t�~Лv�\r�L{�Y:6a���x.�WU�o?�f̩I��K6���z�.K])���BO�b��:�)@�(�	l�G����5����ƣ�� D��/��AX�OW���0N&@$��*ʈ�m���$:�и���P�?"]�g��m��-w���`�=��3�����!�ԃv�Zjr ����]�S���?LȦ���3V��w;=a��ǡͥ"ϋ�����M%�ei�e�RrݺJ�Ѓ�<x���߯�|�����t�E���J��'|�>w��?7�
3��cMS�CL�LܙcgZ�B����͠�n\���tD+s�����n��``K�J�M��$�);!�z���W�5����T��/5�9`�l�]�np���5���͝��J�=�j�B:]}Zq��2����0�ʤ�=dN9(�7��SP�������X�����G^�ѥ�`0Ӷ�(�����<��7��JQ[�4R��j*��UN�⽒k��vd^3KTr%U���<���
�,�Z^	'�C�l=�礂f�h�ky�0�w�ps���2�#�a�=�z�݆]FHi��ȹ��'��bԐ�����&�C
t��[bY
�A('�U�j�+�
H�.�{�PW�`�+�Q�_%�ū�K�!�엚2]i�w��	 j�a��	0��@n�j䟏h7v�����q2��/�k��4NL~0��wBic���Rs_�0��`f���L�Q�6qF�*n�Z���
�L2ܗ�o���r���_-������ˑ3�u4r��r9b��K5W�ܕR��~$?Ek��o��+�P�:���0��0�� N���/����[;=�e[�o-����٤�g�dP�6ܽ�f��w����?)^��ta�H#����8@L�w�R����ʅ"��$�4������� S�Lb}ȏ5=����L,ս��8����1Y�6#)�|��^�_@�rVӢ�#��V���ׅQ��l����Ae̳/)�_�O���㩸�K���	yM]M�.�xX�D���T#����Q��x�����Q<�W0L&^"��ؑT2�OYs��N ���=C�<���J�c�\�箦�;2à�=L�F�����������KJ�fRB��g=��3W����3����µ��+H��v��Y�"N��W��A����U�U6j��n̍�&�: �����d�����䐊�'�a��v�چ�	�鋌$ƻ�n%r��������+5��-��[�=s�w��ۧJT��>�Sסba��o�ʁ҆t��W%Zz=�U�Yi>q�0�%qi(��� Df��]���S�O�W��H��#Oq�ۭ�d�Z��FhIS��~߻��\G	bl+�95�h'�V�� �����s�=@ѵ�x(�i���Яr�IRa�}���r"��Y����E�5	���2Z7HP�f��^���t3'4l����^o��=�	W�s��Àp��<Up$DFl����֤�j������}����CyarOqX|"�׃�!��>�ֺ�����>�r3>)A(8g��4�X�Tϕ������y��_��Y�S��(k�h�o3���������Q s�Z���_���1�`x�'{ut!����f�bʶ (o�
�c=k�:����ǂ�
v��{��SU����\Ds�v.�2.�1�V��,ϼ�,uɌ��1�����K�@�����G���U��>zwŬ��C�]�`��i'v~��,JiUᘎ>(���$O'��
�p���@+�����6�ጏ�C��O�㴡h��,}��hz�UKq�c�KJ��5(�����X�GwU-!-��7qkR�'	vhk�	n&�-R�z�7��Ǆ�<�P!��EXj|���'��*0fC�Y9���3^���%Ud�Dr2�#hv�5��0>>�����<(�V�9b�P�����]�<���g_D�;n��>�S��xy�'ʀ>p�p���˥�A)�k��B�T��7�0D�1&\��g!����$k���'r-L�����T�!h�����d	a��"Y���!�/O*�����9w���h� r[L��u[���o!���+��)�#0|�ϩ��鼶�'n
���c L�����Z��4����I�<}7�q/��xj��	�T-7��52��@��#�E�yY9x*���si&��X��]�?O�몮��^b��anX1���L��x9�k��� �Cyܷ�NѦ1Ґ�~�HOC;X��ۇ�>��+�!�%��g�5���Q?,�����0�c[���R(ɠa�Q�yc$�	���7^�>�5]+׶hv���X`0dx�b��$I�;A����v��b�,	/oؗ�o�̔3�1����V�z ����|���qMF���pו%�5���,o�.Jh�cB���C��d�+p�cgf��Ъ�a�?*��v�*�\����c���S9������E� � 1��x���M��B�4gj6 �c�V�B�+ҕ��b�}<�s��ܽ�׿"�����(�Bh�N�|��[No�2�Ob�1�Mb!T'�eJ��oU78K]���ѱ:�v���`U��X��J��������d+�`3�5Ѷ��u���<y��Vu��j:պia0�;��Gd`{2 G�d씶��O���5�Ӄ��bh����r�Z�l,;��o��l}��ȃ��SU_�PvF
x���7���>��H����㔘�B%�;
��fQ�Қ����0=CArE�R?�A
nX�Rl��'o������s���8��:�*>�z�"���D���zr����"�u���)x��:�v)�1����TAr�[Cb%��j�J�7�4�h�|�lmME�-�EI�NW�z���Cb
>�=?�f�I���N���?��ɏU'�_���ݐ���c������G��*�2������M�P*X&�x�d��*�D��5y�04� ��K�(��FJ@���1;�ޥ��A��4���i�,M�4hЬ�>]�L��N����3�0���~
�4yWz[[[���7v��E
�Y�c*���AL�&�V�������x��Y�RKm�5�Q�(]� �n�z+�Դ؜[x��vn�W�12V���"��/���h:�Y��q�V^��Y�sl[۰F��f^��P���r
iPlk(�[����a�)�s�_��F�8�6R6~�up�BgDǗ)���%��!�*�n��i.0�^e��v{��P��|E��t����'A����j��Ϩ�:5�G�qb�*&N>�e(�B��q����$���xvހ��3�tR�n��[�f�&���Rf��No�eP�GJ�wT���'0�����.e/�`uF�!���Jf]��|�!�`0���bC��]�H�6|f@s����:��"�j�s�p�{�'<){k�=�L���˘�9�3�"-��L�\�TaB�ʰr$j�~���h������Ӹb���s���Yښg����juO�`��A�R,��� #�^h���o�~����GG�Q-f���+(���J�ASmw٢�J{	F��j�����w���U�c�X��9 �u�IV&<��y�P�\ٛ���S�FՍݹ�ػ�VB�c��ɮ̧�-�޵�$@�:b̽�ˉ�83>����f8��ѩ�}
���8�Y�ʋ��,7����"��񡵼/�K|c0,��{������H�'����l��Vne�0��?!�TN�?�_o�=6Y@4��ZyU��U��h�K����8���y��["�"�|��[i>�P��_����&��m�����,%���8YArr����x�_� ��i����$�����7?Ǫ ?R���,Wv��s�-	�r���B�YL�|D���1@�G�iu�|���n#�)[�_�(��,�'�?Yco�k07���0���h�'~:D}�d�;�]�&�f\�w�QQ�W��d����Z�rr�����~��~��l���p�铀JO��ھo~͎x	�h��`t7�uĻ&/Y��-қ�J#FY�p�?Q7�}R�>c��"�݁G2B��4�
D����;	cy�z�������W>
��&Ϊ�{��m�4�$����������N��-�+lf��Zw��܄� �+�@�ݔ�2�2T�t��	��h��O��*��!|��팟����L���)h�}N�`<k>��e
�����pu��'Y*:Hy�}�	���..�fu�E2)�$vN���Կ!><��)�1{��"C���u��Qc���+k%Q�Lزu�p�ML�$HDN#Ku�f5����(��Oz�iT��H��	WO�V%��j<R-(����Y��a��ȉ�x(r�!hq�[��O+.7����5�9�A9N�E�}���H���C������$��5Uj$�Z�>��Dbv=0��u0%B����cm��t}ify8O�c�Ds���闶e��ő�E+��w�2���⩈�z�z�;�ր�:���(��itDO]q��_������PM �#k���_oư;E�)��)��X�����L�2p���j�EVw���#ȸ�=��xH�rQ�~�:��Y	6 	DaXP�ච����$$*�dp��~������J��-ʷ���:��}6�cJH��xw��̌"�P��De����*b�d�;���W.�6�i�~��C/�\qFe�V��]0zby��16��3G�z/"���C?�A�	c���b}�'L���,d��Ď7L�l��3g�|�$-��_3�������yTSJ��aw��ƏT� |/=Pd$��V&��mZ[O/u��^w��=N�3�KZ4n����C�P��9�tC�`�1�5��!�lx�w6=��c7��{X�4U4/n�>|��fY�HH�lz��i�3��3o�@��v?d�<J��j¦9�KRu�wRj��v:�b���Q�^�`�j��$W.�0����	�o�Z�k$A�����ʄ�:�ĒF!c�ý�i�h���`s�y1S�_^��"��
5�
�
`�{	��L���ch)��G�n�Ր����~�[��U���9�Z��;OD�jA��,���K7�铨������"DL�0�7�u�����oEk�\�5{����ޫ]UH��w+N��Ӎf&l�`V�y��*�<L�]��n��h��#j������XR�u���Ʃ�۱RЁ�@ɟh�
��E �[@k��o7;���e�R�`'���R�Y�9�X	�nƙ��,�K<b�r]�<N�H�����CٙfC%�v6��.8�ƉEb-~�*Mih9�H�J��������e�O������'T��� �������,F�x���6��O��w�5�;��vhzY�X�L�C;���v��9������.���1��o���p��0VN�9���)f���BM��,�2z��3���Eo��R�J��ߢu�l��;J�p:U�*�Z��9���Q!�e�V4��8�����[���Z��$��?���M��y��'ؘ���Q�>�L��4ś�U!JL����u�$�>&��=F����}X�""EN����XɸŢ/�7K��0��Dq��S�ovmP��Ab�J���w�~J���8cÉ-?�#4;���[�A�-���E鲨�J�_�bp�w����p����O���'��Z.�T�a����ȁF%������*�ሃ�#DDFŰ�uuf�yff�'ߴ��7��2j��Z��ea$08�T'L�������G�M'�Tq���p�<_���D���\t�l���U�(a�ݘ9=�?��Vҫ��z���Z��ovvïP�wCJD-O`�;�XC��O��T;k8���`,�w���d`�`�~��]�r��O/f;
x��v��7Ӝ-�b��
�yNMz^��/����茷o��",�\(p
Ii�N,��_�F	]/C�̩�Ւ���2�H�>�u(��6\��neF"}���@IO�wCP之!w�_��^]i<�cŷ1���C�yG
�%�
ߗ��jH�����{�#Bpw��Ҟe�k�j�*��\|sKw�u�,��O���<4���V���V���7�{#�V>��D�I�����T��:V揝J�ku)�Fځ�:�ɇ���H
}nA��vxU\��boo���^FH��5>�A��V�_�f��
_�g<8x�Uax��	��|֢�N?x�d�!��Ԍ٩�6��_�v7�*��XH�qh�����v6u����L>� z���q����\���U}u@��f>;{S�	�+����q�&�JY�&��_a����<uY�@�f>ݪ|ek'Se�B�6������ װ��\~�P�^/I��l��|�ǳhsh @{hC5���Ϻ��p��$��p�����K�g�O�4ve#����vk�P�����i>��ƫ����躉��Y1���_���zde����
,#s�qc|Qih�U��)��˿Y�iyl5�3C\����ƙh��c�k�̪�Jc�7�����^ONxl�����ܡU@ȟ�ށ,,��IM��@����j3F� �m���΃�g�
�'�M$�B�V�F��N�G_`0�?q�^��/l��z��4ts�_��o{�~��ѯ�=�e�'7��x~��OWR��tP�BP�8�����T���9�@��v�U�!��}K��;���Sgg�ⷁ�r�du�a���\f��R��T��]�a]��m(4��.9���pX���WEpp�f�����mO�� ��1��;I	s^�a��L�s
*>�m�LY��y6|sI����q�U�|�Ri�뙉K��s�yT���r���	�X1?XB�cpxU�r*j�bT��BR[M8�k�;j�F��ɀ�9�pȭ�bAO{��7¥@,X�է���.���q�TZ�V;������!��(6І\���6�f��ß�!����F����Za�3�+���}��#<w#h#%�M�3�~�l�x���v��uS:&�ue�W&V�ҩ�<��(�n���m�bwG��ʆ�����9�pGݐ!;r��a`}�q�ي��˂�T����߮Sn�eA��JD>wg�������^!���Ԗ��ē�V�D�U�}�!�z���j>h��~��ci�}�i������揞
h>Vfd�>���y-P��A�0��&��Я5=��jU���)����B3��j��W�\�E���Y�兀�Tx�v�3�-Kz_$wͧs7iy�SS��>���)ci෬ˁ3{����Ó'ӡ'��ls���x��1ş6V�g~ctP0��ɡMV"�3�)F�/��pv��/%<ȧ>��p�j}�Qq}��yL�>��p�s����R���`��w��M��� ol���B��c��N�I���z}<�e�ل '���:n(��}';#��|۱=��bm�� ���s���ܞ�݀
O����r �ղ��������k�E�3���Њ���\گ�<��<u�h�;k�u��|e�|�B����љgHy�����4����+p)C�J��6G��|::�W���˞m����Ku� 
H����>�i� !QK�O�o̊5k��Ai��sy�M�{
#��9��E�� �� sB��dh�����9��^wT����)�C�}8���,?o�G��Iι�1A�6v3�}�t�ř�"|�M
i��%�e���e_i�H#+�Zr,8��谇�{����aiLn�0=����}|*��g��1�͗[.s���D�8�Y�Z���.�a�O�ƪ���%0Rj�#�+��|��{0P�y�#�v��<������.���P_����][�i����U�" F9����Sɝ������W�@���s��f5g�/)Ik-q汫WlZux8�Xe+ �3�,�N�}���8�:��]7�^���������rz���U��ߏ�$��y8�@�:�ޟ;N%Fn'C�,�=�U�,�jW�����9�����b���p�/�'Z�Omt���ھi+�Iqׂ�Qs����k7��.A%�t���|:Q���V��.������Bm�l��|�tz������^��KaRP��|���ERO�����q���w�XT�n_��n<�5�9b�9\x����{rZj����
ce��zѕ�`��5�W�"k*K(����|�wJxDy�<|����rr�G�c�6��w+�q4�O{K2��d��2ZY�*��Y���i(���\����ZZ��e�D�3�%R}�7����,�g���+C�EL�.��Y�3*��g���-��d9޷Ϥ3:Lo�g���U'|�G��f��������r�9QDD��`S��9uM�p$��$];��?2C4��Ŧ�VI���E���
Fi��~�G�g�����h�-���XK��c�}&�X��}�a��g�)#��]����p0
�����Z�$[;���+t�O�G�JM邫�.�j��	��16��#�v\�X�:+�D�<���~Jy���R\��?@nC����kJP��n�+q��v�{Yc�ֱ�d󂜈x�����yi���8I�K��]�W���)�w%'��p��m?������K"Hc��ylJ����۴�)�Q�n��Ox?bǜ��7��9�mz�f8pE�ܽ��-��wS|B��Qs�S5�+�^<�0>[l�#$<T>~�;���y��|�!���J${�GM$�Û�M��k�'s�3+x�M�9��$�v��ޱ��%���>_����:��ޡ���kI*kM@�^�q|�ỉ/1m��I[��l�%�O�#q���1v�`�]��!ge�`7�K.j�>��8�CR��l���'�vɖT�������A��ŻP��A�Y�)w+��~��Z����C�C��>y$��a;�be�$���i旭q7��Ճ67��F~�Uw��p""O�V��4~��%��.�i��s�}����E���R`d���poU��* h�V��f b��q��9�MM���mJ��C�O�|m�&5�<�,l�̰��
� �]^������� �H�z�"+Ҩ/Ι=���I���0�FکU7
����bְYu��p�ׅ���P�e��A�iy�?�u�~��"�N~g�輝����і^�9ʹ?�*I"��P#�3��g<�J���f�~��Ƞ�>�q=���k�Y���,�~l���"��ԩ��Q���T�W����.�RR���;B�����M�U��m����� {}��a�7)r��uM�zVHT��d�w��K��c^�m�C�2y����8��G��R�h��@GW��9{~!'���@"�=$VzA���&�\�
j<�����`��K��],�5Q����4��)����� ���Ӑ7�t#I ����!��[`�s�?#&o�]Vo������ư��XqX;� �*�gTЙ�l�~�7^6�<Ӱ����ۛ?���&Ě/ "����cos,�E��'�����h_9�<�*���x ��C�c���M���8maWeC�a�S��UI��+�JS������䭝_r(^3�#��t��I�>4�p�c-��"��F��bb���ເ}�Jx�O��0�7��<�g=�o�P����S�ԔX�}�������q����F�Ҷ��:D�z�$��w�T�����)4�����.3������D�3�L�g�J����`�#�g�����;�P����@����J�.��-Z|��c:��Z��~5;�a2�V��$��rd����T���Y�5V���cJ>Yq��T i�Q��hhT7���YF�2�z�MOOX��W�����e�iy0�Q��^��^Yvnuh�C����r��uL�7� ?�;U@��B��N�Ov@*G�l�L�KZ븖֙s�9~7�b��#4]eJ<e-G�c�Ƞ��ej�͡��!�~�}���N�o���f�"P�w��Ӡ�]Z⣗d2q��n!��4���ھkOws	��xj�wi&�]}Y��l6��'[�_xu��5�y�'��V��l��cO��P�0��y깟�Ύ0�~L��8W�{�w�3��Ei��&��B�Ʒ�w�&%�z�`�����t􆽤W�-�ݮB���Ba������Fqћ���)��bB�hhY�m�^��|s�����nH��eX����n��`��t���ؕ,OD1i�.����o�$[��9�p���x�ڨz���Uo�^v��0muF)�H�A��:NG?��n���xu��jG�l�ق�~I4$�P�����c�۶�>����}��$����qj=�ܵC�ׯEwЎb��M4�z;��`	��;�"����A�x�F��v)��,@em���b%��bk32��fR�3�y/=�q�t�2�0�'���D���<zV�B����c�q�b�MD(k���UoUag�c��a���R�͞S�J�����ޭ��4W8R����.y)�r7A{�TC?m���LrkU%��Vdg�<��	�Vx��>~_�j�y�H
��}�x�MHi��f[Q��6(��:Կ 5�b��C�;�����0���<��G.���Q>;(����2.O�y��"�f8�{)9��G���;<6B��u�U������y��D�@�LΞN՜dG�K�lh��m��J�7W���8��!.���V�&��'h��L�y��g��ޯ�r�юȰ�{���ͅ�����캩�p�dl��
!N�{Z�Ny��i���L������c�U�6?9��aL�7��$��X��"�W]*���PI���PcL���XV�9�n3 ����F�w���6τ3:Qf��O�(�Ԗ�~�z�7)'�����|~#����H������Z�����/w�w�.ʐ��A.c,�Y���'..Y)+sP��^��	�?BKCw�3�gu�Ʌ PM�O;����ص6w�|ޝ�*_ʈVKc��#WeyiHqg�i�굝��޴A1o�8��l�k��!�<�m��(����ruQ�h-��_�S�?�a܈��v��e&�wp91�C�B�K�׮��#5v�Nk6�t�G�hY,����ϵ'�`�۠, ��NiH�"l����ڄ�i2Կ�_�J9: ĠA�z�P�lTん��ܜ��=����N(�$;��̇|�����ݭ���q�UYh��n�{p�I _���巀(���8y�{�_5���̞l-�t�/�<31У�*j�?��Ch�0�/xr %MOhQ�n�ש���.\@��a�e��y؉y�kg󃵥�{mX�R�h=��vJ?��.X^{���xRQ\qC����1m����U�%=�����{�7n�h�bm��;��Nt�h80������eL
�|`�5�~:ҡ�R�ٵ(������S~��Ms�9
���2Ay�|��ԙ�P!�=������5}�4��msl�h�~��ja[4ͶlW�$�.�����J�̎Y]�x��D��^$IfD��'x��xp�Hͧ/l��ӽ�y�|����N�s�J�K�2�./O�;o��.�j��n��
�̓���r�B:/AYMq̻	Y���Os/#:��6d���;,�u����[���/���a�y7@��)���o:j�����yU��/j�R����1:[��;�1�~�Bz�m���wT�|�8��]*k\�n�n��wI�H����ٶ��-}�
O*n�#O(�_PB��":b��8#YGvlv�%ptk�%�Q%d�&�%������؞���IK�w��f�$˲�0�/TN^��۬���g����T��nD9	<=2�ޭ{����~B���o�6��k�V� ;	"��JH���0X[�]�
H>v艭Uʾ����[�u��:a]A��jx��}�\h��+m�����>f3n��;�5���S��o~q�)i?=>�d�d��7l(,}�x�-
�4G:���<YZ�}���V���	�LP����6KF_���ɮ3��;�4���K�E������$���GP��4�;������^+��/�嵓�J�s݅���=�"�����ō���^)�{;X�%��A����]�F1�{�=�wt�!���͜�B�<�_�T<tg>Y��@���.0����u�|���o�3m�	�~�rIf��!�i�%rW�M��ə�3	}��=���L�Q��;y�螒���e�kJ��Ի���M���F�Sa��C������/@�9<��ܣ��O>5�U�a�Y�7Z�U��Z�9G4-�4]�I���M�#+(w�z'�_	��E�����`�sy;��If*��s�����1��l�_��nԮ=k��5j~jo5b�g���ڻ��Z�k��(�j� BIU�Ub�=����_��+y�<I<���9��9��ۇm�KI򣏰 ����fqu��mʍ��6�y޶��H.�.�x^���!XJ��q�I�`��KR	�#��6f�W���~���%�g~�T^���5�����I�r��oʯ������@Ȭ��Վ1�� �f�~���>�����v�e7%#E|���]�C�1*���6v�25N�œ�	X�t��5���٥a�w�>�)��pc�y,Co��J�ϡ1�����*S��;x+�L�5�����DY�ê͏��v�b��7�}�a�	�7ؚ�IK��]Jv�T���e�8w�<�8�?}]�����6�.�Ƽٰ�(}O��"YBy�i�iu��2�/��藨5��v_=�BД�S���</_���[�wgfZ����	\J��q:(���Ҕ��|���l��/���b l�v�?I��$3M���R�M�C
v�tf��� �7�Z��=(�����
�S�rY�4��p-u�RE�KIgN�dmꘜ ��t�*ԋ�"m��(������ 8;0��5���FidVXU{}oċ�Z���I�v�)]��=q���o�p�;���~�&b?.'Sq^��_X���t����׻�=��̓���r�����6.�fu<s$0�_|��usJ[xA͝4{~�pTV��c�K�M��c����u]P@����yd�(������͓Pm�6���`���ư��q�E�9H`�4�HG�|�S�P#�z�$�g�9��$~=I�k��5;����]�' ]��\$���������EAѪ�J"�3��w�n�D���7��zi�\WƎK~Ζ/�h|&�?X-@��s��s���C*n�xY��C��t�]�J��%+���'���;S3�h��ܗ����X��:��Mw�T�qz8����^?�q_�'e��(~?ظ`|����{���a�<\%�T�i�5���cv�f��	��JY*΀a�MI���v+�l~��G�^�����E�|3�/��Z���%]e|�R�}\��1������7���~��笏�� Of�m�so��	�=�+����~L��8.�߆��$�+� /¢5i�^�=�a�����	�7߿Kᕠ	��i�׸��n8���`c���;)e��}�,D�.H�%2�����&�lT�F�+V�$����1G�(��̨����w�n��q1C] ������ޠ�R�R����T���"w��e�W���<۩�"�&��0f>A������n�^N=V����j1�P \p���TQV�Чϑ֭�)�#C����=�pp-��e�M��l�G��kpz�S躩7h}��H]�%M�}<�,�^��V1���Ȧ5��Ƥc�.�G��2������,�}xk�<�����}���%A��Xf̍d�.H��W��oe�e�!�Wp���'�G����ŗ<Am�������;1�e��]�tU���L��."��Q�i����r��P�.y�j��q��x�{'جyJ�.�v�;�O���x5��@@9������kp�ZR}�"�6��Nv���������
d�?２ٸO���:�{����r�aB�^�Xu�p�yw�׫'�"�G�o����\�!��l�D�� 4�>o6�!_��P`��oN�d��n4��n8��5���!����fX0݇j��*0}O��GV�y���ZCׅ:�F�"���ƽ�Ӻ�Ͻ{�z�`�E��.̕�-7�-����7۱'��s�a"�s+�F�\��.t#�tyz�*��V�ɔj��q�-��9�C�<�X�c���+0�JG�I�Zo�ius�Q,��q��Cb=��9��r��R�;��ސ��3�N�
!ra�m- ��q@��(x5x#����{ �!��~���⫟���B����I�b��� �(E �1՗�kmJ����$�(�N0�K���\��)����W�1ڪ���N�z��/2R~v����3��Y�m����0�Ѩ�%�|���i�`'2�9�'/�?_�#�`�_��0�jD� <�'���`���zIHl�o����:��N⏂|~P�H�[�f���d[r�A!�yAx�^�'��� rRn{6��o#[e�\�g��y�1��#j�>��UyۺK���� ��=k���$��,�=�7��2���ϲt�w�a�����3�.uJk��]%Z�V����)&*fH��S�e#�~��N�x��{����x���2���8]�2DX������J�Y�27��v^Ǉ7mД�t�q�\����XO�.x�lb��X�jGyX<��a\����Z�-�i,1*מ[�_���j伂�}o&�rN_.x��l�%��kU0(��,�Iw籫���hӮ���ٌ��B�p_�hx1O9B�MX��\G�-�W���6\�,7<+��$A���&Rl�/�NPz�c�NOwR�Fϻz]n���w�h�L�MXeNe�{��%Z��䩬�S�`��h��T���T.^u�0;�?Sq�Ԣ�3VM!�{-T�{�m���Н��&�iư��R���*3�EdV�f�N?]*��x3�6]�[b�)�Y�p~�I�=4����i����|��=&�2���M)Y�$F_#{a6�@՜ �P��5��w�%�ռM%q��~�M�D�
"i#g�3�\ ���x���n�j�䴭?l����'���XJ�wamB������v�׮ ��B���BꂊD��>k�$s����o�u�+e��c&f~���Q�u���"�B/��t��j�o�@�*�5�*�c�y8|��J�iz�i�\s����7��ջ����y�7�0�Rf@�v��������}�E�F�/ۡp;k$:��F��9݄��9�/H?
���p!ҿ��C^^�f������מ�!�$*�d飷��)r��`'��亃ЊZZI��r9���GMmE������<&��㦶�8(^�o*������[�^���%9���aRL�ݓ�}��WP{q��	рR��� �H�{����q�7���E�O)�u�:8[}��x9E����k�݆�[�7���O���*ɮz��������ޕ�/�?Xg�^&��<�kUdv�9�&�>��A��l�o��V�Ud�%Q����e���E��7��S��
�Ưx���	x��<����?54����M�${K- '{����Jf��h)��ѭ����,�J42c^p;J�v��T�ҫH��]f:�������P?��
�~t��0nJ�+.��ǌ$씄��##���1�U>+c�<f�1�<�L��x�/�z�#yR 7�R���q�/eY���#���,�ٌ=�K[	��)�����}M��v��[n��1Y�L�T�.�݆�=�V�J y��)�[��1<�t ��:����8촆�o�}�p�Jΐ�6 Z������1��>C��S$7�[��2 F�� 9݇B��T�t~Zf�Ӊ�.�s�Zk��'�P��nZ���Ǿ>f���]�VLk��5���*����J�Ƨ�����}i���T`�V���?�CE����_Yi%<i�����+��k�S��u� Ծ�*X���/G[-%�Q���r%Z��ܻ/������د�8��/$���y��! j��
��m�pt�������[�Zp�K]��J��
{z{����0��q���!���m�H��Ϊ��W��\� d�]|i�3�&�Aq!�`=��f��t��a�����IEKd����7��^�${6*��`�ʹ�L������=(�-0=�#K���&����pbb"A��2��o���U���E\������^ʏ�����^��v�YHjn�A��v{�}��R��aɓ�3�o���+�偬?�q��g4b��&�{�uk F�#+���fۿ_�j`���M�	�J�Q���װZ�tS��!�/F��%��=Apl#i,~�� 3��/�=��ص�64=��2�F����ߓr���6��%�X�����c'A��1lȷ�`����J�\\\�e�=tҞR�F�(bO�������`>_.PC�����^ו�̼?t+}4Z���j/���VZ1g��D�Q�W�,�r�=&j�=�Uw��u8H�r�dڢ�G}�@��Mڨ�9_��\?�L�٢k;-�����w~�6���35��� ���z٣��H�OBlb:/��,:���,������1��b-w8*��(u�����Mw�=�v0	Ag��ފl��ʈB�lu����Q�b_����JB��\lvz����f�9c��<]�,��$~=h��SUK#wj�)�g~��W[Q�䩄D�E𞈧إ��e��Ç�^p����<��9��Ϋ;���fh�|�'a\�a(��Q�Zo[F���̦���1�8���I����?aO����1%�tXI��^\̸*TD�QS�ٵ�F��ᗃ"�,�AJ��]g���]�k��.=OU�Q�~A����k^%���������xr�)\���U��q�	S:Qj�Lݓ��J9���B�A�J�\m��
�STi����p�3 Uw�6��s��/���X�C���;8��!.�iAx���-�`�ë�hԭ;�[�,@�HPf��_����G�E��}�+o�����yU㭠_��!d�M�E���o��nC\Z�������%�OF2�%	�F�k���Nn��N٥�c��#�x�HI|�&�1]�s���b�?5+��5�2��&�QY%q<L�!R��x�c�Z]�&mC�;�Fv�k��Ҟ�v����1�8�<���T�_��T�,��nd"k���:f�2�){�]�G�������}�v�9����Ǿ�L]h �{�q�,iϣ�y�h֬<#k�� ��BB1��'V�^gƎ�]��}�����;~�pgC_�~�=�f��f1"9�]�`���v�U�7�)��|��W�N#o�����
/ ���<w�
O���!�X��ٍ)�l�b�IUr��G"$q!AB�<|�pyk��F^�k9����tw�S*���ti�Ck�(���M[i-N�#�͊��R�V�z
W�@�[k���Ϯ���o�)���4A��ߙ�WM�c(��x��Q��/�J�OK����ށ/t��1v�̈����X������j�uߵBr�?@�Bgv�*5K�d����>[��ET�[��7��XX�Ot���/$֝7�#+�Hq��D��n�:r����o���������R��ba6������΢���Vw��psy�z$�AIdā�i+���1i�8g<�����`أv��j62���s��Ĉ����c�¹X���C)&@�`d�@�)`K��!r��c5��7Ϳ{K� ��*J"U`\oD7`��Y�w���}��JH�\|�e�3������}0œ1�/�J0T n5��wBlA`�n�.!j�q��*S��z��<R����{;�ԫ�W^z�8c�G�,�b�r�#��/�	0������~�Ԉ�>��Sg᫯��.���MM���r~a��xg޴?BN��2�s�q=�lWU�0�:Ǭ�����4���'�,�~��g[U�7�g@ Cxw0 � �k�E�$�E�C-rmi���H!MnsO<�[	�nd�U,&ӕZ���C�Vқ�>1�#w�M �I��6�|���ZbQs����7��_3�z�ɱ��~�&D�Eܿ�֣�!0T]���%pG%�(��n���W�B�o�O��|��\�Z�'yb�\,Ik{ĪC9s����u9@�M�iw �@���A�;��gW�K?0o��s%�<�i�	�U���u�A���ϸ��@�@P�����!�{�#I�I=�T��8�L������y�~�o-� 6�������(���S��S�~��S�Ѥ�	6|��5WI�+{���^�9�~o�)A�<&�n~0�$�?���y�j"��_�}�����[��+P�E�ɜIS��t(>�	|����6���� ֜�y����uOX�^DS�x-��^0���a�﫻!�񄮱���}�WH�ɪ+���564�ֽ/��K5�7ԝ�4,fUW/��=����g|ĥ��L���f�<�z��6�y7C<?< �����@LQ��&�@.��魕pPC[>�,N6N[�;7{e��7K( ����o-F*n"�F��R[���∇~T6�ܮ5kQ�$�1]��2H���4���ϑt��h�
?m�������%�-�9����jf�;���74t�׷[�2�WS|+N�O�����t16����[��
�S�+'ߍ�K��{�vS�zj��!�-��1���4l�q��=��8�G��uu����B=�;5!��Xs�mEc���ƙV�!�r7��,�s���1�A��0X 1�Κ��6�e� ��Ժ��,U�p3�f����##��>k}R{�C�^�O�?<%ЭlZ{�BBqj}:��5�J-���lk#{,.���� :�B�o�(>��!	,�i=�TT6=��9�\r�py].�HJ-�Z[5���E�-�O��:?k��R-�i�H�~],<���yqf���~(��ړ��P�,��������&�����r���t��������E���a��Ѥ� jd�;������&^��`ڿ��
�8��`B�L���8<���B�]�Ģ�ҧ{�]|W���ilS]��MX[����&6�5}��zr�@�%��oX�;\UY��>��e��YT����n��tBn2W�*����P�+3 k#��*�񨪑aGɦ7l���v&���-g�?ۂ񽺪��	}E���P㩻������zg�$��\�DLW��H�z�qѰ� �=wHid���1I���_#Ij�jC!(�$��L�s�\���8��mj��˾u�*L�*
��]��Ө�RWU5�d\a�3a�Y��� �S�ț��n,���~��3g�k�6�������%%-�I��M>�!�QES� ����S>_"g�
���HO����h,�h�C���5	�gBݿ�������{C�F*t�a���N\�u��ʓP��H�ҾL��G�����λs���DB¦�կ6L�:�`�KE�h����hj���`����W`�%�<���(9�L�~�=3���C�Q�� ~S�)��ǂ��񐭂�y
���ݫY�����l���@�v��h>w�#1��?��j�:�u��ެ�p� ���<|�'X�a(�1<7����S��j�i�;Պ�d(�:������6�LP��}�פ�ִ�3��r�6����K#��l�&��}����SO0?�،�֖!8�r��p������m #��3��r�ݗ�',sq���/��TIQ��O�S{��G�4~S��|$�%�fr����@��A�nf�n�����xmvG����!�Õ�)�j[��<�v0�aPtq�NY��X B����)�F�o�w��/0����fr��\hx��F�q��kl<l���{n\ap�#�\�#4=�,�w�+��4�
��Y�+j��?��6N�E�̀�	�X_��Qw2�s�R�v.�Y��7}�0p��Ƨ�����t�P�msYId�f�l���������U"�=�l�����g�	��n�k�����a�z�c�O�L5Ds� *�(6)u'�>�`�����n�4]~�*[�9-G�~P��S�؀��tHn�o��K�N���B�� �)�R;�q���[�'o�>�-Zf���j��/��[���X"N�ח�y�,]P�$x�b���
��(��כ�5�%݌��?��P�~�����D��'i¥����T!^�:����,U����H*e"�ω7�w웅
���S8���"1��*>�>H<A������/��<���n9���ż�kj"^����}�D���j��9��㭆29b}{�;>�elc
]�L0�P��} ��FR�)��Cv�pg���U���"������>�H�hT:�i<�n�wŝ� �o�h��e6F�|h���55oк}7l���?b��Iv������j�bɅ�h��l��n�Ϸ�y\����^�RFLXz���> $~VHc�{�R����H���@�Hm�5�4š##��f�w+��f��������94�nh	td�b�U
�a�8�S)��|�0�3�$����Wcڜ߼�2ߟp��#���&�J|���(j#V��N�]
D���4l��yTs���Q[�a��~�p���}L��'M�����k5��;� �h}|{p��M��(P��c�I�kA��Q4�!� SNSx�����Oڇ�MW��F��m�l�\E�_���&��|~�K��5'���E� ��˫M`G����*����%z�q�|Q=��f���<{������K�h�����84�^�L����h��-�q!ʇ`�N�>��^�v:�\2L�����7:�8���Q�ؐa
p��0�J4W�O"��bW\l:��������3�t����}��;�"�E�]��"H��ocV�˛���g��o�����8\ԋ�Ȧ��	F=Z��о��ZRn�Sk�t�9	�t�TL�<	���e/�Pd�>&Lj+�0������F Y�}��/�J>vu��~�~suus�az�b��|�U^^X�/gP��^��ay5/E���Y�xqU�FpQ�?����>�=t���ܓһ�Y��ر�ȝt��3�����W�r0���s�&B2֣�x�F�mb�k�Y�5o#�TD�gDuk��_'[b#`�0��}gӠ"\�ۿEӁ5�˳�{���u����Ӓy�"�\��>}gO{S�d��ӛB����^��[Z_?�n,ˬ&�_����SU��J��m��h�S��G1�,J�c~���;]�w\Y��}}���%�ŋ���TBK�x�x�^���yM��r�:@0G��K��+�X�C�p��m��H���t���>�!b��v��}�2�-(i��l���"
\d8G�ÙIO�92�?�LI��9���{#>#��[ؙC�Wz�ѯ���k��r�- x����◸�����������q�=�A�"?��S��`T����{1�X��&��������֮���{�@(���Hx�$�A� L*QI�ݩ���}a�v�N�EZ+ԋ�7<�.LP�BV���cql"n�Z[�\v� �7�i�>p���y��v�������6=>��%fGn�K�2�.[����>{b��\MD����G%�h�'J��#8L���=W�+|��X����mt�`ʴMԪ���;MZ8�� �ŝ��W���t�ᓛ�������:����R�X����M�Tǒ����z�F �c.��`V�FO��Ck�.��{7���w(�3���a�}�4�B5E�n5�a�z�Xe5u��EԬ�VR7��Z��G�F3�rp�_�����N�@�{��6�O�f����[���S�H��T�RX�sqz;��D	V܉��mi, g	�����\�߮R������E���wz.�H���N���������y2?�9b7��(u�1�_�KM號=M0�a�~�8���0'��3��xT]���$�\�^��<�($�͙�5kx0wm�ɾ���*�<Hޡ�����w����C�p�cyd"+�pgj?{J���e��wU��'�)�(��
G^��*�9)2�bH�]���7�@��4�bc��B!OST=��$X� �f�G۶�1��l�X"O�#N�\Dw������P����!
%��A��'yF*HТ֖ �[x��`|�<�2�B*0�lk�)�7�ʪ���-��&� fx��@_l!O��`��a�0�+���{X$μ<�,�;}@��(T�JF�YI
���u��Z��759�^HF��Qˀa��i����{�㠸XG����\�'wr��-Dp�+����0���,�pn�q��V�B�l�^Qv�^�]eh�r;|R嶠�X����ݦ���k�"9��E��[�q��-Pꩇ��h-���rZ�&Qv��y�k��	��Orl!V9j8H�/�6��{��3wO3�M���wK��D�Y���O�;o)\��.:����D5�4S<{;�y�h�Zg;߽a�O)�H�pPt�y�4�Y�wf%�bȓ�7+�Y_��#�m��QW��B��BM���nkdj�"̊�b���qS[br�)�CA#�Eb�D;��C#ܶqM�����)9�Ѵa9�Rͪƌc��H��_q^���܃�'8f��yv�.�D����H1��M){�dwz|���;����zC�K����,�V�TB�ar.��	�%Mm���[����@ZqwJ��K����y����A�d��/@�����T�������`X���PWF1'K_]��;�����V1q.AѮ��+�b+�`+�������ѱ:���M��A!" vყ�}F���"������%�AL��[���sU�FdW˖���[��|jjj	~Ƹ� l�x4��r5$n��;�U]n�l���v�.�V�uِ�$�{�f�0��	��g�'r��e0S��KFEy�*Bimuu+�O��A"λ^q�l��D}�gW~[�w �؍� �P��M�/5;�u"$Q���<L�T~J�N�$oo�#�O�����b���Cb�`5 �SH��:<�m�vJu(�ڞ��Gu��ߔ�4r�ݺN�&Zm��̌ � ����,���ț�X�������?+������P*�@��t�]�G��i�m
L�v�׿�d�/c��P����������w��&K
�f~������
�k6���������󑂷P�BW���G�t�,E?ah�"++����Z��0� ����P���v)�k�Oc2�ޤX�Rp��%���w��eq���0�3x�xD�x���%��J�u2���O�����������u���b��9�r��L��O_v;R��Q���&�oi4oA�zu�~}�����݄����^��4x��l{.}��1�䫎��5
�����0���FCi�;���D��
~x^i��O.琛+�����I=�+pe�<�i��=����a� xq�1���.�0R��i��_��
�v ���u���7�!`mn�i������������k���`�\x���|ӈ	|m��K�����vr )��J���M�Tg�L�	��M�*�n/����.����k���G���լ�X"nM�X����pG��O}�$:!�R��\4F�)�y^\�o�Ro�aDa�p��D�&��R�l����$kkj�\KgO()���#�����W�=�'�c.�<���t	ɷ����i�Un�SC1�����`�ռ�\f(��������&��]��5�oA�y]*o��.{�� M�I���~SjR��C6��B45,y���k�P[����+�qlCp��fOq�}�*yR�l�%�̺8��şNrP��*>�f��+�ٕ�:�d��9��/?�|��d�#C�ߴ�i��2C��v7��Rq�����#7��8̘���c� �p�eI�[�N\��~�w�Oo�}���Wn -d7� 4)���[�Nl,:�V�Nb�m']�[^ �4;�G\����<��{�8g��::~���tR�Y� 3��K4���d���
(�x��kg/t��pU]M�]�xQ�E��)6��z�>#N����gv�ɻKfǣ�{�5
6�+�V#�ٖ���$�㗭L����؇~�n��j̸�����mq� g�&�^��2��Cx�f��G�{�� %���%cZ.oq�)U}�83 ��R���tQ[]]����1�ȸc�҂��Á�m0�~������v�,�O����PvK���wާ����������#�5n��
7,N�Sa�\B����D};���.Y �����l��^d�ήY�\cSVC"� �S�~��'��	?��=U����O�e����s���%c��ȡ/aXrm�-g F<�n)$��p��.��$߲���@aq��|K�٭0��.ƾ�>K�1N\�����\~�`l�����4���\(�O�X|ڰ�ӑ� ��r�=�� �i����.�z���6��)���GN��/o��-�]���,�?��Ͻ4ă�
{�>�'QLy��X���Kc��-�e��sFU�t��4����{&(P�)[�KP@�v[2Ȳ�ɡ�A3�4��]�q���Ⴟξ��ʓ$}�D�����~��,��zD��j��z���ӟE���'r�0FV�'JS��G��&"�F�b�BM�ܞmF��V�c� [(�P�w�SZE�9j�,���r"IM�Go�Vt 尖���})�;����t��QEM��8�zN �ˤ�e����.b��̬� ��UΡW�����I핏Wd522�It��a�uMu��9�um<s(�7t���v����:��nꔊ@�|�2�qh�Y��L���D�OdA2��V���Rc�9",�!�R�Pį���iX`z�3���oqYC�(uf!`�)�O��j]]@pȟ'�n��%������,�Jci$��5MM#j���^#�>���eV�Q‗�h��y���HL��FY"՘_r���] ��Ҏ��6@�XwI�߯HY���k�Ï����j�2�cզqN\�ɉr�.���pT��~4L����WLp���������+���6��K<���\�O%%pP#�EO-`~q��e�5`�`l�짪�u�I�E��?��[Lq��F��x6� Ÿ�p��摷�2�3�	h#>bb��𭦀��?h�k�WL/�Yt�T�E���]>(�q�`�/�����=u)��Qۯn���g��6T2�5�b	]H���Fp�L�ˎ��ȱϰ�8X�Ks!Ao5�$^[�ƓQ�?��-�/�uNWϿ��T$n�����#�����뤉K���l�{�U͠�r+�O+���$����D�,;��y���L��s˧�[`i��&6�L27��Y&"���~�(C�yy�=�޿O�
Sr�\6j�D��]BGIB�E����#�H��L�@v�՝v��$q+���j�G+F3�G?�5�3_u�9��(�EM>���џ)��/W�~!�%�/�2T���xB?�`�Nd���߆�J �
�x�5�- �m0t��[����32t�,�P|�)�sC�2S��
� `gPeTɐ��Q�(y��3��'o��fԋ<<<2��f?[�k.�(7��6��-��%��t�����Ӷ���������߿�J�Ck��~�5X;O�8�����e-&{��}&'�A�)�(�����v���ڷuc�#L��Ŝ��������
�?�/�&�3pJ�N._I|9zԃ��}��`��^'�J�luwu�<!����X&g°=�w�m�:��f2�X���@�+�E�̲k�翹�hO�W3��y?R�˓����w��b���d[p=#$����l�oP��UyI	��6���0�Mʳ�߶h���D%vG]����U�$}�vPD��Q��2��e�K)�p��̆�����uL�62������''�.Ve@��s�L��࠽�Zj�f�zbb���]��_oeVb�8��mK�h��H����XA*��b���7�e�z'߁�2�����u�k};$b��[	��7x-���ybW���g���u�X�ɛ%֪��o�x�߲}{@y��4�N��?�J>ȸ�Q&;��ûa��v^�j�m�)4�/Ǎܠ�Ü�f�bcKò�|Q�!��H���nnV���C�(R����T�PfV��7Ք��4ESU�:L��"jU~���	B���{i�%Be�)��J.�ZY���=ܺř����kaG��P��3�	�V_@C?�6m��g|���w=p�ܱ����ʓ.��`���� >C�S���?6��,���,��^�� ��pZ	���b�J P���Wȅ>e�8��)��e�	��JH\��9��H=G(����b�/6��D����m���}3Z,7�
(NWR� �����r*��i��>%��~/�pG3hx�.T��ڿ+�~�;w�}����<I����Qg�x���v�As���s6ъ@h{û���"2ʥZ��MC�������3���G���ɀ��-UM���Ǜ6�j�ֈ�Q�Ci�E�Imq�l�XE%` ��]�wM�J$�>��?�E�~L[���`̋�������֋��YH+�4 ҁ���5���������(\��P�r6��� �r���5(W���۔��O� ��7@p��|�Vi-�QQ]�1�q3�;P�&�������SND���D�2v0h�:(������hR�<y�cu��p�t&���ͤ:�ڕ�&�ܧ���]b�䮁��i�]\����G_Q�h���S�o����>EI�Y �y�f��ٕ�Z�c4�������9P��b�;,��'π"�
_H#O��͚��T�e��0�:Փ��r�b��n������J��ϩ7Ct�ز�E˨0*FnsZ���r����fSTn�j6�����J������8�u��xg^
Ӊ�Y��1?�tl�@#..'�k�f����U����c���*���)z~]�������a���,��=�B���ݫdԋk.�k�����@'��`�C�?�m�U�Z���аT&E�W�ۯ�-�\Y�����2�+�J1~��V����-�gk�R��yyy�H��hQ��p  ���\�Ía�.�Iep���,���,lQ����S��e��Co(����&-�`n0��}��R�Q�X�6L��`�o��\A�Uf�Y݃e�_v�o/@�4��ɷ��~�4�7!�<	�A3��X:1gۣ�k�
�]�$R��������	~1����%�] ����%W|�����ٶo4PIq�m�%�E�����9�(�m��f �,�� �pw��+����9c�b��89q*�9��rS�2A��p�jފ����d7�Y�ދ��U�?��T|�>��~}�F��c<��Q���L���V���9߹j�%<�c�_�{v����&�t+z��Y�֯���o����΋�':&�[����'ԩ�~�T&����n)�,a�8����?���!��`��ۋ����R0fȮ��
wp��ܽN���[��J��m��ơS84V�t������3���-��3Y��A� N�K�k;h�~���<E�j���lǉ����u۝*P���=�>#�fZ�~Q&w>2�0oֵ�ã#^) !H�r���%[��c�N��|��o�I���� _C����*Sl��)nAW�߂n��?"o��J&�"��w�P�2|_�Ď��t/�E�/jR��%$S]]R\|k�� ���g���?� &^����߄{�z�5^}�����u\�d�.�{,�rMj�Sl�}��c�����Np����'��IZ`�Å�%��1�|�Bh�T����b}0'y�$�v���h�ys}1��Ǐu�o�����a���N%���d_�R��ԁ���|�$#�FgR��C1w�;�{oS�̋"���p�b[�0�U@;�E2�|��?b\�.��@�[E�i<�?wj*RAc���?�ӱ
6
���;&�@��
V"V��>�I��j�F�;��8�$�o��w���3&��)���d�]���W/�e����H$n�i�+@�~v;U�E����QbL}��x�e����������nǓ���Y)�#uC�.m����X��,�
u�!��k&1 ����#��,�9��[�<<�/x7�O/"//�ah��(�M߿=���Zn,t�Q�������CBN��UB?eI=�/LN�ozj�b�t�h}a��J��s��G�8e��w�4hQRD��hP�T�2p$u��������jKՀ��fͶ.L�>�s��m/�f�Q�c�?���Waø��?�����X\	��.���R��������F�i-N����xȘM�1.���Xc�-�X�C;�"dpأ'�ò���|Z�P����ǯ\`p�FY�I:4L��\Ͼ2��{ڵ�&Ԟ�n�VWL��^Wi���U�����͐r��E+����%�R���u�v��B�g���fsÄ��F�&�`}��R��@�Hō��3E|v�>Sr�=����#܎����4@��[s��Tɍ?�B���p�c��v���:n���>�C���fT�mH�p�b»�^]	0�񀐊W���6�x�Tq��r0�U�����G��Ey��vaU}J��j�kL����Q����/hk$��� R���߳�뙴(�Z$#��;f� 2�N���f�E	�1���O.���,C'�j�}��&n�V���ۨ���i��ߟ_�SJ:9O@ �$޹�E�|�ŀ�n�x" br �sV��\��$�?e���n��8�pDT{���*{=x��(nn	Ȣ��mZ��]�o�x���FV�t�v���|E5����W����! �0M�^0��w�ct+� �O��$�E���/���[�$��}9�������Oc4�l`�ŀyv �5�RP��[�g�8�`��ǚ�2�ֺ��g��h�wt�E'~�[=ʃ�~6$���$�����G���A5�=�Ž�[G~[���2S�D�Ȏ8i ���N���3e�K!��$D6��A�	�l� W�&��������Y�c2�	O�e��kU������|{v��:I�!$Cf�5s��*�N�z"J��Ĳ�Ѽ9�<�@�ҷ����Ɣy�� }V��`0�6���Cd���&�"Rh�08�'տ�  b����@21N�F8�45L#��:�Nf�S���=���_�x��?wiA.���[ (����]e�_ε�d�md�u��g>9��{NM�������u�6��E��->�:u� J��1f��H�������_R�d���d&��.�g�+!+3n��Dv�^���uq��y]#��J��������G�۽�}y�s^��8����|��ni�����M�_	��~o�y0�!v�:���]��0�tH����k���˟6�� ��M2P>;gT��<��C4�Q�A��P�� @��1X����Ew �1nD�W 6й����3�)���������+Louq����@���Ϳ�����+��0n;nuE�A�<��_���MoJ0C ^�Z����Jbz���Պ���Ɗ�W��ή�!.4t��ÛS�X�]��`	��o�ǔ���;]:,U�V�{�J+
L�+*���tݩ+x�+���_wQ�.�:dO�R�]��8�<*Q���-ܼ'���}ì�3�gb���*?VRz��|�_Ww�:汝4\�`��#�JH_����{9���m"N,���z`cp�*��,�=A����e�sG�f�}+b��;�|���1�5�o%%J��AU�L���	�R�Q�x�u;�W���� ��ț�BjU��0CK��!����P�J��g�k�}�SCo���:M3�=�.y2��_�6�>��#�ȟ]�s�d�ߛ�\��@I��g��C��]�pSk����Ů�������pw��[d�~�PA�C�� �e��ת��_�	,)��~�G�]t���������5٫������~�Xφ�d��f�
�@	�"�O`����?������n�ǧ{R�ߦXY���SY�����~������՜�_?���p���i׳�>�������#Ns�7��U���&��� ��7�����]�|*P;��,��"�]�w���y	��J��*^>���R�X����".8_7f䫒ϋ������
����-�qL�W���|��P�|P)�b�W�L����,G�d���zb�P��ږ��$NsI6���)��tKh��3�V�=�����F^�_cXj'f�ʒ�&?��h�mk�@w���,���{/_��!
�7�l9��2�7 P�gf�y&��A}�؝}7(�[�$@������A����a��B��5}�|3C�tJ"��ɋ����3��]���orV����Uٔm��A�Kx�&�x�'E���~M"�����#f�f]R;D?i��U���xhg޸q�$B���s��s�#.ѼA��t����dxh�n�}d5��{Ƈa.�}C�]�7�l�T��<�	XT��
t�8?{�o���";UaUqz���ML�?�W��R�3�"
�n�7)r�ӏIp�'k�S]����!�4�=L��q4�� ���y�y�����}���gj�֍������!gd ��
��?�T2���7w�����Pέ�QKgFs�ԇ/��݇�n�"x�v�w��G�m�������cA:�Y�Ԏ�(��Y�N���gײ���Q# *	��(�%����C�M#F��m ����?i�vaE��Mvˇ��j5�����H���7thŠƵŞ��T���T�C��� �7nRq��$|�n�'Q����*�ض�(|��]��q�J�1m�S�*�d^�� $m�ͩ��,�e?¿{�:�2l���#O�&@��ʤ�Z@�$\���nDEѧ��0keV-{�%۬û�o���|�Q��U:2�B?�v��yS���b�=D���~�Psq�P0	�}y]Q��"�fP�A��a����%n���t��L�
�lj&�̹�

�u�3σA�6��o9�40���Z�lߙ>,���{x���a�L��TRu��F�m$��c2��ECC �0�9 ���i;�����ͽ���\ߏS�'����9�E�`�dr:���(���oЊ��Y��{n��)<%���	�{{z�} @���T��'��?XUY|�Y�Ǜ3�>��~�l���K��(f�����H�i
�]��+_�E�v�m_����T p������Zz��*D�R�vviV��q�.M�n������W��9��õ �"7�ce�k���rǾ�)u��|3A�tf���r8��J�F��L�e�!�6�{W���؎�ǂ�{��bUr��4�9 �1�xh!����G��lB�ٗ�PV�..��r!���n�*��X�+���
?�Jp�d�� N������f�/,K���.��f�����\\S���7����T�����s^ݣ�=�ZDZZav�m�,��Y~��S-{�/�a�f-Cf�-�W롶��na��o�����B�:Q���N#Y @Ƕ];��gY�H$���AڬW���!a��Q��e.�B|pȗ���y���<���K���3E�;-��N�i=��E#0^ёX�l>�7+��ao�9ģn(��pS���U�8R��)�Z�����?%В>qy���]Q�:�X-�Y���з�c����z�����G���{h���u�ę�G��tx	}��|��(�/�?�}wZ\���m�
ƑQL#�R�l{���=$�O�qK��О��;9o�y��Qn���Q^�t��DH�3����J�0�m�ۂm�1�|����_��5�R�PG����"���=�=�������Ұ�|�a[@35��#�A�����ުO�C�Ðp���z��\Rh��mz˦�dϾ�(rcF��s{�h�#7��\��Q����y~�7+�.k9����P1ʟ���o�j�׫)9�WJ�X���?�?�S�]�7���/f�|���w.�'O��u�p_QT���&�L�����c�y�:���Xy�F�M,������荇3�D��W��I>����iv>=��_/H+��yc�}��Է]|�p�����/&�|�ԙn{g�ʐ*�J�<�8F����n�HE�q�JH����Šg�Amb'X�'!S�	-�������?M8TY�y��=4do���/���^Z�og�#Pu�O����E�zYmj��ʓqE�	5D�"'�A�H�Ot�8����(K�*2�8��|=�-i}q~fp� �`Ԫ�9�eyS�b���{
FCb�Ѧ��	��=V�\���k�N�˓��Q_�
�&a�Gꢷ;�������:)�����ﰒ�.������|��n���)���ެ�q/!��3Q~���/��W���$?�ȠJ�hh@��$vRl���t���}�J%�:E��t��B�|1&�a�'k�R"8n9!�W��R=�*���S�ua�>�+!�&���^]Ơ�9��8�7z���[9f�[_5t[�;|EZ���ҷ�5K6��]�/�4�@b���(�y]F�`Րc�9�@�Q�n]��c�8qԣѭ.óR��a�q�ߚJ�L���م��~w��J=9�GV��c�4Ls�	��h��xƏ���OPOަ�8�p�7�K�3��<�}:�p�Z8s�!�V��q;�H�
ަ��<c6����[~���� ���V��c���#)fTn�x_î����t'N���}9<������P�d�z7�e
��k��n����ޫ2P��X^%���*��7i��+�Q�T᧐#Eլ`y����P*[�� ΑG���⟽́qZcɡof�7�SM5����c��o��ǘz�s`0�Y�>f�:�����m"#\�=L+�&��l��5�Vj����ʚ������}cU�oό�a�υ*J<a(��5MXy;��h������~��4êS�عwsʚۯ���&�G�����|t%���.9�F��44O�00�N��R��H��Kq&�ɗ)�q��a29�I5� Î5�IM�)���H�bS ��*qX~��C�6xM�/p��j�V'p�����-�;-1�"y�dS~�Z%���$rv�[�I�@�*%	Q���	2���ě���~ic�f�C>R��>�կ���LsP�P���}��n�BqW+��d_Q'a}�TN�n��ƨ/$C��C�b�xФ�j>�=�_DB�#`~j&�Ψ��F�g�X�_�7a	�]�v�/���{ݡ|����Z��*6 �H(6 ��������-LrrrC�4�4��a����Xޓ:�	�4�n��{t�axK�ڕ�c/u��DF;è������o���$DaJ�d|��_������ː�L����-��c�R�V��b���&&!g"�1����ߠ7�.e�����Y :�!�:�M�(�[I/t��y L�>�����[`19�y� �/q���q�(9�; ~�۴o0���r 3oq(�qk��gSVK�_v�}a~�����J}t����j`}	g̞I�y�8���P���J[�{t�H��'���9Q�!���E�Pk�����v�F��鏆��V5]	�G����pK�xʄ^��Q9!����C���?��_��;)���xB�#UT�ˤ�p�%���7Or�N�;pb00�G�y.H�_E�s�Pp%���a��u�G�� �:�j=�z�����^VV�n����1V5��׆��f���Z��*O�_�X�w;�J�g��Ci����}O��FG�CtMG��bS�.*A6�e���/��Q�����V*��J�eT���b��[Ӯ�߃� �5c�}u}iIx��=�z����3>ڭ���j/�wC4=\$��w�do�o"hf�6�a}'����c�m ��t��������R�^´7
�?��T�<��[��\�XiH�22�K���2�D�o-��ts�Uݜd}2!V��(.F$`m*I��H�MQ��!!
�g���S�TB�f�%�A���v\��c��6�ҕ��^#|lH�>.ɘ�&J���:�07��Yr���i�>�$������ (����e�
{;dFW�T��j�qqv8��Y����:�5�|؛��7����5�gC���sƈ�^֊����ݣ�z�k�6�_~�����UK�,.%�w�� ���U�8:�S�z�w��!�L:EF��#���#�0�]%�!��2���ܬVF:gDde�}+�5�督�	 r���1o��z���q ��?��ٽ�YQÙ�hO��j�m���O���NVA�dDa�C��Ɩ�D}DkY������=n[.G��r�It�Ԡܖ~�̣�k�U�q&~V�+ؓ^�5A�� X ��lv�o�~H;x�6+�|}SE�$��3�S�b���F̺�"�d�dBy��K8�g�fr2y��[wqn���|��m�V���&�2�"�������[�06�'��W�k@�FҘS:/�e�H��f99k窿���ƣ�������TXܼ�>jJ[`���T��|�/����m �<�M*D�Ƽ�rv�J��/�����,�v$�f���N�z%Nr*h�))��^9�$�(9�c�P�p�:��ש���㞫_F�5�<�;%g��e�{mHi��MT�S���		��/.V|J��z�މ1fSp��cg���������0�A�;��<�M����;��I���l�4��iV�3 v��J�{a�e¥oN�I}3kh��Cť�l���^e�=�y�vk��9]Q��.D��a��L�����v¹�u(�+e2�U���&��<4�N�%��o�Ѭpg[���L��fu<N�,�4�w0%��a��"�W3%�{���w�}Cq����vA<	ӑ<��z3-׆U���R��Zr�S$��^��o3Udx�xݞ�����>�d������rB}S
�me��L��8F�
��f�ٖ ����ᝇ�"J��@��#�դ�u���?����n}���T7��;X���Xl8O�?Jp3�k���儚�"�<�3А�����y�Gn�Ӄ�N𸖶���Xu���iC��oEؘ�ϥ���-T�H���V�~�!&�^��yW��J�z,��IY��B��-��K��S#c�xL/�aKN��s��7�@�'��9��f���a��`�XR�J���<�/.?��"��Ar�eS�?[z	�99���p�{ф�#Ħ�`��>3Ʃ��oR�jy��D�ơ�K $2B������3���5���}!�{����t8������)��!ύ��?�3��P�� Л�r-/��z������ wV��Δ$s������y&wqP�Z5�ye���/�:8��˟Ύ��iqww�LO�ц}���	'b�$�	��ɴ�1����y����÷_H
@��?��[jz_�3ұ{�X)�-%A�� '�$��5��0��I�����5�::p&Ü޿��C'�U�i�NV������% 9b��,D��u��~+�ֻGd9�[buvC����i�Q�oޛ��q �f
t�0`��k���I�q)� ��t\��ޗ�r/2m��7J^�z1��[�:�w(k �gݙ��o�R��"L蝏5������pP�� �$О��!MOJF0�H��˂��I0r�y���*��_R%���?��L�}���L�pB�ř����I�)l	\����6w��!�t-N��.Ɣ[��	g�2l;	o�r�Qe�%ab�[bO~p��B�<;uѳ"���2��xq��بl��,���7�+����~���K�(_��x
/����!mV���%�(2�>�eXG���fT�lP�_�%�nꁻ��Y�Z�P��?r�s��]5ǈ)���i��{WFLEB$�D����Y����:3Xh���R�Y�I��.�JYF>-���[��m����qP�~�oNI@x�7�zN7�*ԩy��V>��z���Ez�A%MSBo��#�w��#X���*A���m��.���a�׆�����4�"�,S;���ջ3��������d=Ȱ
���h�X�ٛњD&u��'�h	=6N��k�K���:���4�&���1N�V����H�RL�>
��z{+�����_�(o�i�c->�1��F�y����o�(��@���8u���-��=���ϛ�-�x����v��F�q����p�L�t���Ec��<���zz��i�I06�#��a���m��	p�9r����fS�ukR }��T�e��J��<L��V_z!ˇ_�dfZқ�Y� �#�un�ॎR��o�o6�_.o�Sa�ɫmuR�L|�o?�98�'M�z����<�������|��FՌ��҅1/�:�H�й���O"�/g��c���+�Q4������ �a��&�+Z1��ز�2�~��c�ƀ�����5)�C�ՠe�����莈��㚅P:	��;N��Ds(��Q�\e���;���_�d�u*��JW?��c�G;�/w8�4X�/��U�ov�Q��r�� �������D�;_�f�w�_<t r}����{j���V�z��t�$�#|���,V3b��sxw^���ڟ:�4U~U���'�����?�u�K�Q_[��<"�?�"^�?�����u5����/��d�����r�H�vj��?g�\ǩ��˭�YѡԘ�nu�;��H�J�v:���K�?�j�ٗ��*w`�=�ӹC�����wQ�#�<��ti[�xx����%CL�����h4R>�̼.c�������+'���_:���O� �y���5�>å��1����C�Dsk����-�KM�WC"��|�v5;�M�e�Q�� �(]�E�����#�^���,44�j>s�йKG��Ƶ�.����VJ=��a:�z�iE�1O�6yPI� Xw�R��a���m�KW2�a'�J�i)cu�e����J��J�E{P/�R�Vg�}8}Í)vsgBZ˞�r(�sX,H�I;�7^oO�^��V�����7$D�=T�Jd�rk�"��g��ω��$��๯������B���n��q�%�Hm��ᤧ9]������h����y�������Nt1S�2)���%D�;T�%T����~u�F��i�}�
��v]�v:�G���K���I��]T4&���{_���	��2`����qD_��6�9"U��[���i�����2M��ۂL�M&���@�V��N����@��}�a�\��/�r�C�����6�g�Q�s]�{d�,�I���x-(��L�!4�ZoD��<Jdyι��햒R�A�m�3aIބ���U���|��>)���xc))�s���QY���U�:����z�G�ĵ���<�3k�J�1�Pql#�-){)t�:/���f�({e`$��6|@�fH�j������S|��`;}��f�S�`��"��i�}+_tsIÎ	 ����j'�g�3�H5��IۧHroO$]��[b�_N�g5<}�3cT�J�����w��?�n?گ�K�������96?Q"\E��(j��Å%��Ẍ́C!	xbb]Pq8���������+W������'�T�=�)�bU�Q�B4)�oA�v�h�����ib�$����oE��ŋǒڹ���;qMr�������=�_'~��8��w��m�
N�(����H����lҷ15�MNo�ȭ,ed�R�P�&T�ӝVv���4
�g�n �&���1�S�����R�Y��DV
>7F/ѫ���Ar`���(#�Zl���z���@Ô������a�q80M*�>�����0XB�vGj�C�3����nvC��N����'��'�g�'��)I�&��.�gJ��M�;��}|�[�uD�����,�=��&^�FܘbN����#2���m��B6�)����3���sd;�R�[������G��*K�g97�O�6�f�����#�yf80�O^�8��v@�!0���,���6�L��- >M��Gp�0"�MG?c�{�TxHE�I� I#e��^�����MvX��:h�KBFT6��d��vɘY�?��Pr!��+K��~�_nO蟭��E�����_&�Y؛p�I����?��t�=�)X�.N�.������wS+eyC�B���� ��	S��Y�N���6����Ҝ��KO����T �qǡ��?�����a"�0�
���_h�|5�/�7�H�q��Gkx�a5�C�����}�1�0Sj'" ����G�2�$�vx�\�R&�%E�L!׊u���I���w��Ͷ/�&���s�jjY�����/�5�"`��woXR�9+2v���C��<U$��t	�+/�咰5)�Y� F��&����x>�� XNm��4!䐚)�yz������D��:�mɻC�@��!�Y��t@�m���#1.�G�-�X%%��>U�����Q�>m�����ie��}�ר���+��G�+ҞV�}egON�����2Hr���Ws�����K�v;���y��0���} o�.m��,�9���b�FFZ뿵�G�
ѷ��ƽ����!��r-����Ԓ��GT�lk�U8g�h���U�z��iIoQZq%ڥ���&4Mu�]�Y�j,35�Dp��|^�J�ܤMu�}��K�y���a���2I{�1�%�,�s��nN����%M��$ǧ3]�[%�x%*?�:�*��X�LÖP.�>���X��oD���9���.�ًj������2'L���V�t�Q��-�|VNH�.�l��YG�Hx��3���b��a�9��߃����o�؀�OMp��-#H�d����}f�?_� q�M �mlo�*���J��(����>+��䥫��z�ݼ9i����_AAA�����H�ʇ�+���W=�P���(���G=^�&/�*A3OV\BkF�d�+�F>�V`�M:���W &���`!��^���Ҙ��(��?���H��?�%�i��[��O��������#�y�\�&�X�	|w�|x7�M�"p�D��=Ԋ-#������l��Ցc����!�K<�Pt!$�x��~�ng���9�ź���v�ra?��}�]��=Zzw4� ok�A餌(A�e-7߰�ڽ�`�C���b]"�#`^,׉�#/]��j&�9%B,.�@��^�4}�25����o�r�����I3���c~xM����Fm����߉kw*ݒw.o�Ad�!<��,N���~��-gw��]Ȫ����#_����ƻ��$T�~��[8�3�+:��Y����T���j����[o�E�7����v�@��t��o
��ǨS���k5��%3�%Jz�鏋+�r�dڅ�*����z���r $Μ�0}L�G�d�b����(�
 k؁J�&�~5r ��Ngu�qc�X���N��^��Y���]�G�{hEw�s����ޝ��h�i+���5 j��(�x;�bQ� z#/2�\4��pp��Z�3K
yNX]���+��������ᕞ�Tgw'��D%'�T;�O�)��j�0[��Cn�O�K'o��h�M�����P�+$����`�*�����.P�.�9�~dLػKO/%�њ<�<Dl"I69�kS8b�`%�F~�o�#�y"�O�0��g��!� 㗞Y9�vlu��SR�����}k��>�=\Y�ᠬ��K<J�:!o��_�t���L�o���`�u�7�|C'�2���L��
a�*�����)x*U����M��>�0g@M&�7SIUk�T�������!%_�V�Q.��A��h�hO�NL������v��M���Ӿ�����v�﯊=�4�b�7g�M"׊�խ�P���`�����LUu���N�������2��r!�ˇ��?-`��<��C��o���������h��7�;)�Й�ZZ�-w��V�/��.���<���i��,54s��؀Aҵ4�]� t����� ���n�S$B�sR�F�^�������8|�/�3<୘�y����}�?Ad����#�>�ս%ܰJ��4;�{߶%��eO���u���L��I3>XC���`�ܮ�lҁ9��H�^?Ք��;�x�'֑[��O�����!K{����}�uH�Lw���n��42�wi�o&���a��ܜ�sj���m����nrN��=��HYlmd[ˊ3�v��Df-7��ۆ*G��w[;l��A=U��+��Z�L7Ef]L��
�ǐDv��]-=�tt�{���w������ބ��t%�h�gH��34�������	>l\4��nc��!1)EU��0g�ܴ����b�7'%����ܟz�B�δ�d1���*-��7:/�'�N��Go�3<�'��^
��a]d'����r����Yj���ר�$�`"C$���
X�g��[wҗ.����$�yN�v.��nuK{�ո)�T��(t� �~���(�* �`�Ą�`�TU�m [����L
�|����D����T�m��[��,���m�A&�Տ�Z�и�������x#�շ�+� ��#�uFJ�v?�
D���N��:�`H*{d��ٽ��-y�Z���ϖĿ�1�<�������-�WW\��$D�(���u��H��_oΊQ��z���?otڙ+\^�L_)�������1y�SVv1��
>�x�jJh}�o�K!cy
�G?�t�G+?�L�F��N>����X�З��~~�ܱ{?w���$  u�����p�Ν�Ε�;�$zQd�"z��T$D��6)^O$�C�iJ��~�'z���W)�P��RETځ ��7�ر,B��.?�������B�1ݜ��C��|��t]�����W(�����F������"�u��h���f�t
���#~^$o�������b$W44,V����hz?z<��H�;�}eو�=���^�%��8�0��F�J2�<i@�w~��J��eF��l�}Vp��g�z4��h$���E�\��uX�i��.K�![�����9v�hf҆��P�>���������+.�_����Eoa�8Օ'����Z3�L��*/G`^�������`��*�ߪ�~�,��Ŏhj����_��;n�B�FJ�;����3e�3=��k�,��"�%�py�s\6ԭD1�~�S;���,���:M��oz):��(B��p�1�p}]��_�wC�>'��n�1�K�>��Z�Z�@����1�ɞ�gKl}���3~��2�dv2L�]1�W�4/���|�G9큸���M�3:�&.,�#���f�iNJ1�,����x��7���l+�;ʄ�V���n����iδ�t�35u�%��T�d'Z�&�%iʓ=�JH�"ʒ�K+���@B}lQm9���!M����e�>⋋���2Y��5��'����-���y6K�@���&���	~��0[g�^mIp_�,��o�Σ����}�2v��F\�QLR�I��.�jWR���������@��p�r+p�Nz�g�Wߪ�{�� �ѻH�U��\3�P?�y�e��햱��a9�:�g�|�jO�oGp� $9d����>�aq5i|�7~PK��~� b�'�~��73�I`��ު�Q393^3�ݺhU'��Ҩ���0p)�%�z�؏��m?7 �P������t��B|�N����>fxr?�:'����^ͭ�Cr�KE-�-�s�t� �>߂�E��KQ��機c�y��2���P���(�Iܓp�OZqJn���A��!���[���A��E�/e�|��U4U�V�ۍ�����)P]�!�6
��0z��=_�ߴ�� �͂CZ��\2��Q��?�� �Ϲ��,�7��P�%ة�>�'���i��Ьf,օ���J�5	�RO�`������i��
�
�@іE2I�ޑ�4�,(�"�l�704�?9�X�^t���T�?��s��m)�Pa�Wֻc&�Y˯Q�kVf�^���ȥD���R�fu><��"[�V�?�(ߟ�K5���A<H����fg�f^�i_:���-x�iBk7�=R/�����%3_���пo_ن~�ٰ�����+�vq_J��o?J���Q�q��Ww|˧	;1����/�(iH�<p�Vg�F����f��������$�X_1n=�;?ξ`*.��_ �&�KE���"D�M��mŵ����&z�� @f>0���^���ITK����'jr����!�QΡS��N'�z6�4Eϐ�-�w|�!�`���3���ځ6`��6��N�h�d�W���^;�`
�{L@"�����a�K��w���=�v����>�v������d���q�k����и��,1!٧H;���n}�쳁�7��H�^�3ӲVY/W��!స;���o��j�F�ȯ���CVU���1y������%1k��,�����0�xz����	1 ӐN�Ij�I<����9^�R��/�D�cId=|eX��ڴʤj�Y���W`��܅ű~X��"�S�}� &�k���U��
<�M��{!�Ѥ�r��x�6����}[������ xfӷ�Rʇ�ҕ��r�����r�2N�Ob�X�]y:ѿ�c�g�l�y�����������
/2SR�hE�p�d���᷎��0㝇�U	������~������	��T�cߍ�H
`�6:<��yL���CIs�|)���q�����{�����
YO�t�c�(����f���� � �`�����oS������UdH���I�h<�+ӗ2��t|�l��!���#=ׂ���K+bX|��@;V�&}R��9R�ݬ��'>������5`&#rmk0>�o�Ʋ��s��"��,|��'�7T�X�[�	�ZC#��sm��z")B��,<�$���=B�Di�|b��8C2�`��W���c�U�i)�j�A�����JaJ	Ee&�}�'"�	F�+�����&��
>�Kj:	�����*A��w��& ɤ�;o���1ᕻ�r'3e�c4�g�^��0|����i⮅װx g{�ĮC���L{�x�o�6��l,��R�\�� ��Oc+��n��K�#�06���"kT��ƃ��v���]JUѐ�����@�������˽��9X��C;���~��騖��dߺ�0<4��`���f��T��KΤ�����	�Cȥ ����<fK���:�kθ_�2�(��rS�t m`ˣ�?2!8�7p��x�`�P����a�V�������H#W>�9^�<��0cv�B�8�Z�z/�6ݢ�&cD�Pc��e�v��A�<�����)�������3���ozC�)t�x�),ǁ�0����j�9����ي2����2��57+�/6����XN7zVd�'�X�J��Vvd�W�w�)�z���o���p�X�\���(F������:�A�����;��j>���=��]&u�����q;dU���j t���G����*m�o��0��d�播�P��B>�8X���0;:Ӓ�E�mN�1���h�������������3>�4k!�NV�����<b��vs|}7I<�e~��_W�𦴇mn���(����a��X]s�Q�np����=6�M_�@���?`���`w��)�W��	�bbrl	hN,IY�W�����Z�j/�����#��ŎCa�&Bn��0����@d�:66�]���V�C������kNnn'�%X�� ��k�U_����t�vu]�)%E�+P �G�_�ގU�8��U\�$ �n�Vm��=ԓ�w���ꬠ�fU=WA�FU�@�,����0��w�B�{����S������ˬ�6����ZQ�t���N�ǋ=�v9R�/+B�՗��p���!�W��5��T�	}X�pu�˻w���4gS�����(B^:��	?2�i9=��xK���7�Tss�v2���]��½0/+�lW��󕆊��2�u�,'�/�����_���3�ʏ����Q�č}���?-�[��3�rrr�B�.ӾSb�G0� }��[G�^v!�&�6�޾a�bs���w�� �3W�!٠������Vi�C�������ܚ}R���_����rN� U>�V�"7:�Om֒ON���I_�:\8�����9��?�������)kx�1����O�,��{{k��+c��^-N�V5�����oN�j���������|W�t/m�佢�ϯ���)��ɦA������T �ɚz��}�.ښ��0�Ή��}�
@��7�*A���Ak��K��S0��aBR{,#�_k�PM�Ջ;>�(dy������ϳ'��^�|�<��&��������,����p�5��C�srMank�j���A�����mB�;�&�h?�����ѿ��C���
��)o�������펑oh~�2H+];eS������� ���&�!��լ.�J�w�� �?t��f%�Ѣ�)Y�9w�w�7�u���ks� O�<,<��v��I�����w�m����!��p���Xכ�S5'�o5��PKUw��u��\;�&O��/�t׉�PoـJ�6�~�+��aနTBy�b[Z�� _�׆�U>`�|d<Q/E���xL�ԸS�(�)紐�1Ы ؔ��]�;&��!��L���&a��JțNh���b�˥������C�Eڠ��"ۚN����(2f�&)0,�P���B��W=߷~&��u��/VI��e���B�tC�R$F�u�����{2�M)��uG����q>@&�j=v��v?$�_�9���G�Ҍ�O�q�"9ti�'UO@��{��{"�d�>�����2ux4=hj8�|M��ù�1$ϾO��6��X+�@gF�3
r
_�t��{~�vtqѪ�E���%������c���d=�2r��Q�u����Q1g�J�j!��O���JV�dt�Zb9I7x�M��Y��s�����:�6)j����3eu�G�i�W|��C�AE> �����	�.G�CGN�W�4e/3�e�m9u0�<�)������C����}uPo�y�!�X�L20�EN~� ��� =k&�M�!��b)�ɂ�#h`�����o����V,K�'(�?tk�7څד�L�ȱ�����t��/��o��Ȼ���G�9��`C/~kl�$a`.椇��Ծ�-t��z��lò����U�7�⹌�PKġ���ύ�ʘ���c,�~2��*�9m-�.V�A\It,~�'������29!h28x_�*˃��}V�V�1Hv�ϤDJ�S��Y�)��_�R�P��8T��8�$����ce��.F\��=x�9�Or6�n��{3k�?�Z�e�_]�!�������L�8��=0Gv\k�Y��N��{�"��N|J��=dl���F}���g4�����7�3#"l<-�R���7���NF,jY|��?�ײ'�B��,ɂ'��/G,�����~�w%����!���_��J F)(%Y���nV���YIGl�U���%gi�m#W�`�nHܶs��]Qsl
���;���_ѕ�q��"c�+�;H�sb�|��{����Sp�q Z�z.}������&o�T�T6(�ʩ>%i:<�p̨�D��>���y츞��ݰxXe�OY��xbu����i��e$Ϳ�����)��~�H���C���pW�����Q��l�q�+���o�W8�dz�=�T�:>�x����~�����
���#/�K�rS$�����.����G=!,.��Ǚ�1�6?�B�,I٦��Z2���"��&�rs�f<�W�kqaI����t�L{� *"������3����3��e�އW���^�L��t�#;��*-8��s�D�A��M])ʝ�+?���`�^�O�~��W��x�6�r{���!G�ڼ��MU��.�!�|�}��?8�mF�ާ�'��W�QO�^�t�X��B�댆��plv�w)��`�u"%ս�g��U%>R�
Ǣ��U׹P��_�.�#�g�U�%i�����:7˄X�]|����[�~FoS�R�6r��z2:6�B��S�%*8��ĝ7�(]놗���N?<Q�=�N'�tz� R�}�bѾ���,���h�ڗ�"�@X1�B頽�dE�A�P9z}�m�+�`�i��Iܳ��~�Z(t��N0\��g^�ߞș�vq'Rp�:ď��"fO��'v��N����hoD�b�C�r�H���HG|y��_���-���e�����.�FN{�.�S_�E�>�z��5ݶ��w���%��O���恤�A���d��̆cH|�t�^k��J�+`S=�2�pV~vN���+��4K�V�d�+�[Lj�cUO���ϸ�{�����k)��K_��Ɓ�2H����[�D��S)�+�¶`w&��]��������� k�{�@PA�7�*M����Bo"% UzQA��� *M�tH�"5�H�H���N����w���!�&Y��sf����{2����Ss�3��n��X���{tT���}�5�eV�}
����k<���ρ�B�s����<r}�O�{�*E��;�f'y7�*��o�/w�!lI��h⭱"��������J���Ҍ�g�Woj5�[J�=mv?����1b��E�J�����]7��Oi�����DH=#X����Aڈ2���K�&F��w�h
�3��l^J唬N����U,�=��#AfZ�Y̾�+?9����i��r��M:E?Al}�PgI� >U���9߲��B�I!��~� ����y���+������^�a��C�J���B^UTT�"��BR /�Y���p
�JWt�4"�ocSz���b��_����(o�>��ԋ)/�Y�7���ۂ�] $C�0�p.���:�}\�:sZ�n��\�^�rn �g}Q�'A���;�ƴ8{�^MP�$��%h�V&b&q�̛}T8TCC]]r0����㶴�
����%�&?�x��a�K����Y���������d��Q^a_�	�2�M8�-���i���;wZmj�&!B �M��cɷ���\3�_���0D�X:���\`蕗�ϬI�\	���i"g�T~���C�Rz�v_�'��
0}re���$���p�ؠ��Ѣ�&�Ĥ��H1|�9_��� \P�*"G�^�6�X����EԺ����߸r����4hx��5)]RE�<��*{�x߳��fE�8���Cl�W=ҳ�c�y�/�s<��h���=��k4%��kYj��m�m��#�r����E7���v<�6j�J)��I 
˨s�9>�t�L����
�u��锚�x� F��M�P�� ���H�v/�b�� TV�bhѱ�Ҹ��"�v4�[=O�Y��2u_:+P�?��5u�o��x�Ue���&jS��B�Yi�b�Ͽ�����&�LE:������+��j����O�Ը;rǐ�~,n���Q%|�59�愺�Pإk}LPh�u��*�xr�w>�˰�v��vq�e�@V>��y^Q�����<`Y4������N��V��)o��Oh�r����\��]����g'pP��41y�\Z�[롟� 'w8�{����,� G�-� ɌT�p~ %�߸�C��O���8�|	��}�=��?xv��#���>B��Ws��-��+�	k��Y��	��!�髩��Up�Y�o-�i���� fk/��S�β�U��������f�2Β��y@�A�d�Be�s�+��%��CР���o:��Ċ_3��{�ī_AMw�t�U��N9jV��]���،f�x��)=><x=�F�2�|Y~�S���K������bڂ���Z��fo���k�r֩`��R�N�4W{wؕ�*^?��Rқ�PdT�Z�8g϶7��LVңt)��!��
S�Ŭr�Ju9��u���?�9�d�g �\(���xW����]��\�4��C�!�w�$։Ïk�����ƕλ�9�鐬%���Ȋ���
������t�	f��D��\���ISK��.=}��R��Nk���Ǘ��y&�Fǣ�S����{�at+}�-</�&,�Z����pZy�קG�%�����4n��I����y�g��pܪ���'�E��:�9؝��D���U�������:�nsKW�V����b�q�y�_��� �(������B���qi�?8}_��4�M��"�p��0�A쨹F�1\`,��⭎�Ac��ߒ�8r	F�"OG����y��b��o'a�?X�K�ۤ���Y�A�gs�;>u�[�(z���yNj����p�(�l�͑�wD��A�?O��T��c��]�e�Q� "�� �CNr��`��r�ݽ��J�O�C�M��}T]�+x�)��{l������X�>�G�/�|��`� �9�EbX��݂�y=���#�G��K��^�	&dg�)�Yv��]��i��x�Smh�����<W�=�O��NS'97 �|d�UO��JL.ڕ�ƒ�.EE��U��xlUVQ�z�"� �g���(��-���V����|��&������X�!5�	���qvQ������b������;���c޹��g����h�|g�JF�����RL&�ۈ{c�u��uu����L��
�p�����mj��Iv1��G�ǽ0z(&���~��q�U��DKk��EJ{x���zP�]�°��v��BVv�']�pAF�U}F�*#�4*SҸ��n�Y�g��EL ������-���a��z�`����.~� ���1�d�;}':r �1EV�	�$��T]�5�(��I�Fe��a%�V��Y␼+��f� �El���t��0��q�p�x핾����-�Ƀ���B��c��'"���}!J!7��D��ݣ�a�L�vf���]V~��G<(ox��N�N|I�A�8�/�'���drJ"0!H���"bW�р�v��O[����b�d�z��M�z��U���:����0}��}r�|���؞V�x���o.�C*ѳ?0�7�=��1�x�J ���3% cgd��m0}��CO��u���>W��� N�}��R&�$�@���o.�q}O���U[������;�z�^�����z�	����`�<��⋈�H�a�_9����.�i�m�V�1XB�*
�<o!����`s�}���w�/��V��F~�����)w����1��w�(?�	^���<��ѧ�-X�gN��]�%�Ϧ0��˴�Զ ,��ˈ2�Ɂ�6�� m�漾(Ὢ˯ �8U�k7�p�ywև��K�U�my�A���Z�nw�gnnn2��m����"k$�
��e:�K�E��}R
��b�񨘛�"�)����J�I�\lܼ0O�z�����m(�\� �{�U �+�oX�����xf��e_W�/�ͳ�E}���:�M�;�Ĵ{�/�f�
��H��a6�v��T[� �;��l�զ��P� ���,2
����j�.{�0��l$d����;f�ϓ��I��ټ�W�#�W�Q�4�8�]�/Y&��r��Gs��c��S�o��㆝{ӝ�"�~�C�sKe�*�>A�$�+}�vp;D ���0(���k0�Ȩ�w-���=.\��\['��^�It�O�,��Þ}z�ߘO1�r?���,*b�W1W ��c�'��	G��)p�L����u��ofj[�i�m�/ǋ��uё�͛�R�21R#���g�cz��Yn��&�j�=�=�a�E��qx19V���,s��	>��=� ���[�kW���^�k�U2�'FѼ��n�����km�?+'��1$����GTzT5.	�9����v7� ���F��g�Y�BD��������ǷSo�*�A$銊k[2䫱��yeH]����X �7O�����˒ y�駸��\�'q����V؛$|7�l�ۖ�F�����$�-��Kz�*���"�Q)>TTT�Z��_�ng�l��Cw��=� ���ԍ]'9����|��2r�+�ɳ��!����V�*�ݷ�w>���LD�����=��n����^��Q���V�"^۾~�"�"M�K�Uh�f;���	��j�P"*�97�.s���r������p��k��L��pɰ���jה����6)��j���oYڜo���� �������i=S�g�.� ��L�i��B�3lWWY��xi\�LA�1x�������O���=�e����]<�t �Pd��s?�K��Ze2]���*O6�!��'�m\���m�?��&��}�������P*;��U�GD����}/��o�N�����=i׎��}���-�GȷSB�wGʀ`S�H���昮�l��6l3-�qe/����͑��I��z�tm�%KnP���
�sJӧ'$��}��S%i=�*Rs���Ywr !>ؔ�.R��nt\q��󎁖bi��[c�Ғ��F�\��7ߖFG�&�۶&H�����@,~�Qk��?R%;p�Z�����g������rV0Tb۔��KoU~-ה��ûHա�7�~v�Ϭ�Mvd#E��= ;�5V��Z�(���G�W�������{��{�⮿8�.���?�(�Rw�R�Z��[،��tZs͝G>�Ǘ_�n>:|����H�_t��M��B�n�eG}����1�Rąh��V�E{�~�dݢ.�wU�>�֜Q�''~���0�wۡX����`�]�=|���ܻ��y��_����D+��u?��P���\5_����$~x�kk��y��άBZ�Fe*��m�B�Mi�6�HE��[	�:O����0��N�c�}e�a4�g^lg�z�3������q���n�����&�訩O�nS5�j�f��mpE{YG���IG�vw<B�z/N�>:4�c�f>K���S�vX�sZ��HD����3S�[K�}�@,��4����9��5g���w�͡/���� .�l���p�<d�V-pFM^}�{���d����j5�Dc����е�5ٚ���wc=�����|�ߎq^�g�;����c,�I��>���R�5��CL/�'>���m������2c����̦�̲���X������nwj.F�+���k��3��FX�N�Wm�Z�_�"xlUz���*D2O���.��%64Ԭ��\[��<�"4gHV�$��w3�/����#����d�TC����~%v7ӟ���3���*�ʃ�3q.�HN^�DZUȔg.�ik\m
�LP��9yH�q��j*GJ��;��g+�|�)�G-��A�k-U�E/N,�+�oU���,���N��9e?X<�|12�Cb�t�N�e�lb8�w>�W�U��7鶾�J	A0|h��O�><���Xb�Y?�5�V�b	��wR	�g�a���*뻥�^��d��}/)1
Y�ԧ >N����|!���gBH7?<�M�ל�-��m<��M9��FJ���/iN�g4�?"Ñwp\��_�S%�>=���:�@���Jn��B`���1_n~(%<X��-���|lͨ� ��H��^�]����B:��L�I}�zvm�S��WaA����S٭�/j`�4��ǶND�.�����D��Ow��̗�i� �ă�:L*{a��>(��
Q�v*�����=���k>S�y�.���( x7V���>˼ꈊu�<�j9���)z�C(���as���ۯ�Y�$�S�*�t>��xx�f�����M���?�R���{�"I� �4ԔOY?8r�T'	��82�\���{���\���}����w�r��c�"�����q���l2!�S�t�듟���͂���7ۂO�%b��Ғ��>�ώQ]^���WXT���g��J��f:$������-M��	���R��`��[r^��t�Z*U�$U�wb�?�	K}�X%�+���u�	�2�a��Iڂ�Ϩ.�|�#�w��fْ�_l���d�����67��|��Ż��w�P!+��|�k�j�t+�y�O+�`Rj�U#���mf]�֢]�`���}A��ÐK�~�m^W��_�7~����˕�]4��$;����(C.$>�[X�A�;���S�lҞ����������c�c-f)�Rg��ot���I1��7��@2�h�>�'@����^��2��8o��sqf
��~T�.dJG���p�Alt>iDGMF�(� ����9vo�W��Hh��␶?��SIQ�d'y-LQ5oMh�"�O��=�l4X����%�V�S�[ޑ�[/�0�� ���ρ>�?G��ͫ������
߇-�)y�gx+L��=[��J��,��w�4�wS���,�|�ї⤾l��&��*���D��^�N� �^*����d����2���c{ץQ<�&��P�C�g�ت�]�s��4�`� �?噿���Ƙ�&�~u�z��d���<l��$���?��'���_)��2�C���`}xn�i�������s�.8����B�Aʊn��><u�v�����Q^!I�Q�F�Ӳ �(sH�+W���[éƚ�e�J$�"�� ���Ag3:PujC��Ѿ �)յ*���a�B���Λ7�K�ȖJ�Ϭ��X��ᚹnFl4�&D9�{���G��7פ��D�i]�+�~�W �L� 6����R �p��C��z�Qsv<=�� � B5r���4�]�*q.Nv�5J�hj���B�i�ǝ�m(%	��g��|����Y2��.#�6�){�Y@f:?t��1]��'E����I�p��ݍ>~\O?��ي`L��׫�ΊV�֨��O9��Z�]�;�t����:��J��	����x:�����a�T���[��n->��{vԂCs�M�ƽе���7��W|{@�T�^a+:V�.���r9�@ULך���{��;!��X+I��FR��Ã=%�|��%�L6_դ��5�1A��e0�����{������^g���������]�^���0y%���A0J��7o��������f��5YύΤ�D�9���`e����e��i;�����0�C��	Hk&U:����Fѳ�����~��9eRE	�����Y�e��P>Y5���L���&��OC_�uq�x0�V����KC�ȩ ���~|��+�e����\1n�'gd:��}:���_�wv�)���o7% �S^A����,� ��
�§E�jy�|ױ�@i���Z&ac�'�x�ѷ*W��:�*W��$��q�����eA�^'���7��J�Ѕ�'�+wj\�C52T-�xm�	qt��8�rR��5����]�µ��,u<o�̑h�H�Q?���'bE��[z1����}ĆE�C�)X�Ch�{c6�}ine{k�V�=��1�Vn1ahb�w�☣B�t����l��I�k1�]H���BxiN\5�Ca�/��)Q]��_z��L�e:�x��9eqn7�ƹ6!�A%+��fI,5��8gʖ� `�F�.{t"��{���P�WZ�k�g�@�'a����K_����7��������)����|�E�ût9�n�.b��Z�#�܋$��;{t��BF�<&��-!�����k�,�wN���w�|�)�N �N���>���Wº2����ei�s�}.��!5s��c����=��
)��,�����a~+���m����ID�j+��$�,t	~��%�\�4}��]m����Ri�W�����	��w����F�$�펤<�8S8�N��<q�1�[��5c��o#�]�[�� ���v?Y_�r�~�+lԢ�0�%Pym�]���j�yu��V���A�y�F�W��^���PzS��<rW��dlp�����@�"z���ǣ�u�b:���O���ƣ#�~��*���r�����ߨ�/���.C#U���F*Ű���VN�gҹ���|���>����h�?��z��O�[M���HKrժ�J����WkF?<��v��e�I{���'��FO����.��$�7+Ҳ�\Z�yo�P���C�A���+���,�}� .�i����k���8�,1�Fa��q�iu{w��X�D�ڛ����LW�v��)O��˼�$��bך�_%%�������y��ҟ����[��ӾZ7�-�'SX'=�����U(��9�\�LTĶ������՛I��^�D?(�@jEq�E��,(>Iz�
V�*�y��W͔�v� ���v_T¶�#��`~����������S(�Zmǖ�����I7�:����UR�S&��)�������}&����,=�{����dqP����݋���KL-ӏ�ĝ`6�����+���:�"�h+D�3����E�2BnWv���NKz��ݥ�[�M8i�B�ג��4���G�3F��xd�V*��10�U�=������Y��H��o
p�'��E��L��ɏ%��qF�1�fj�WԔ�Q�;\p���2�?1\�"������q�8˕�����3�`T��b�*3[c��5��R���a��(���U}���]�M��#�]5||l^�nV���u��'l�Q����h�O�'����J���o �/��)$�-}���Ѽ�o_��k�~M��.�1�	]~�p<j�4��������)��#�9d��k|}yTLj�6���/�}ޏ��b��z�dS�1��;#�O\��A��[ N��e�� �Y�B-�(&	�y|���.5� �ca�p�|^V�� .~.�`��2�qn�9�T�_�Ŭ�R�,qBmJ�*�
��{cE�I�H�=ӿ�¨�ư��ݜ��{�Ҹ�{�Kg�u�#+�V�����9|)h9�J�!"�2R�o:GS�1��d�:�vX��W��eA�)���d�zu�Db��տ�X��A9���jJCN.�|ܙ<
��D���?��V�{w[�`R_�t�ZoGBx��	'�����\�n�m���]�T��%���7�<1����΁�E�?���r���;3����G����g�w|:�bS��O[�:��A�?�7X .�ŧwy�.��ה@]�YX�M��;�P���V?��:ː�{� �r���͈�ʃ�Խ�������⋶�&���_�o�o�&��>�(p�T�����݈��/���]k��y5�נZ��I�}��(�_Ĝ�60�0S�+�'�����ti)����%��z�M��E�f7��\�u�����kb��:�y��=q�b#�t?{o�<��z��U��4��+�u�Y�t�|�r�l̓c�wj|j|��o��D311�d�yZnb���t���j�H-4@ {���m�i�	���W�=0Ťd���R�����k�\�tf+Y"X[�1����uಎU㭋\Q|�����a�׿��]��S�M�#66^�2�P����b(���_w(��=�N�lb�}t����h��th�۫-J������8�فӆ˰���*����|H��";l?����f'{�v{�F���`�0�M/I�k�U�%ҝ ��Yt71Z� �D���B����������� =����`��e7X��Y�R�i��k�nx�!4̢�^�8�Ɵd�ȉ�w��Yf���]��Xߎ�T WIL,e�(N"\d.@��C2.2�;�Uy�=*��m�)��J�p��|^Q�"���D;�a&D��6��ɵVr��fN٢>�����ӝ��e0�P��o��u74̩!lrė;Y� �J=$s��;kϔ&3�x�碻�/ 8�/��P� �$�JPg���ey|^������%#R-�>�a+�JraL�Γ�d����|�fk���C�o�9T�t��B�	�c��R�W����!�,�͍����ԕ�ᓼ�Ѯ=��,-h=D5�>�>d��8��z���&1z��6D��4ݒN�='�?�&i������(3OW�/D{d��2�<�=��"�6���g ���7�(^?������:g�F����7��I�}&*/�4Xw����.�W���g0��3�%q��r�V��ڙY��r���˳;eQBo��S9^"
J���fY�����Ҝ�|��"^^���cBl�{8�Lट��k/%p���s�����xMkr�^��*�s!�Q�Ћ�iJ��Xv��wSui~������X"�@���W��was_���Ӕ)+�ؖ��9���vWN�=-f٨��|ɦ��$Z�^:"���o嶰��,���tX�����?������I��pwR��Ƒ�t��o���WE��!���3嘐K������^/�氬M#�
I��5-�ˤ���fa�P�%�q8?5��?����@��$$Ҟ�Y��o�aO��Ӟ!#�#���0�vʁ��w��V�:WٱbX�)����>~��]S�踹�^���L\�aH�����}�17�ɀz�V�-`�4do����^�f�Z�d˞��S"��!�˭��y}�*'�Q-7`�;�ONW����Z'�_�n�1��ho}J.�Y{̢y�(�t?���L��-�B��Jwk��z�-G���,lo%a�q����f������VE�R�$���m%�%�ϥ[/�vw��z���D"�+=��&Tۺ;��(��lJu��<�[�ć��=f�|z�Agm�j�m�)�E2�˃���8yϭd�'O]`�p�j�����p�.j��e��m�ظ�.��hL�;`�P/�yV�9�G�P<lf�G��0qN]�.'\��H^�)0A�)�)%�w��A���z�顑�)X�$z��7*a`xҟ��/�Q_5'X_�'7&+�c�dZ=]�f�.[��k�������见x��N��~���-K�7�I?���vb�!�/V�~H���\;6MD��� ��������ӳ�k��
�6-U;�5S]�҆.)���Iί���T�geKզ���〳o����b�*]y�>rJ�
;V����#�bz=o���	�1[�n�L�\z��waD����덤����%̵���Ew��O+�ew	�h'n<�C./ll��*�ϣ�Nj �oVϽ���$�^�j�W
��tL:���\w,�X	~7���	@(G�O��v�*/?�P�Dͥ��M�ݟd}u\�����~�Q��6L�bS�2Wn�&����P�;�jsp�S:3�&4cTa�Kaj����f��X%-�F:]dO�
 1ޔ  �^
9�j����w�ߛ���a��;+QP��*�A�+8��`���K|�āEK�!�nn�����}�����Ml��=jeߔ���\/�j~���4 ��q�|-]�d��Q̕����a	f������xm��ھҟ{��L�NܟVB��ޝ;����F�e�"��n�ʜ��Iq��ݭ��ܩ{��#�ŕP�L-��	K�M\�⽗'��wo��-����d��c���m�L�{�<Aߏb���˝JRz��ćW��V#l���ؗ}цN%L���Ɇ,i�!�����ꝕ<hAϸ��sU� .a�j�	�`tW�%qp���J�F�ݍ4� `�t ��/�������G�/��nlW��:���>�i�b�9%t����_L�Y�LaW��Jx�Ö0&5�P��I_�7P ��D�:v-����V~K��۴�W͌a�z�c|��V�Ѿ���9)�\ش� 	�3*��bd�(����(�by��f�AD{��m{«#��E�l�C�~`������읥�29�r�1�B��cØap����r��/�ȏ�0��j���}m�mU�\q��=�+��#[U��8LP�gr*�ǟ*&�i-�9��
\�<Z�O��;��B�|.�.xuL��mn���g��P�s�l����|�uzh��
I��,�чn��%/��u��~!V���R�$����S_q���V�Զ���"��\�9���w�r�����j޸��+?|��#�4Nko������@��r+6��:�{��a�K��i�- �(�/`��O7���e�{��/�>Ӽ~�l$��1��4
�t;JѼS��o��ȳ���d>c�N�`s����?���YL$g,�m�^g�3�je՗�o�>{����L�Oֿ�]G|�'�-���	p�i�4���
1���D��pjUiB��TլU �H���e�P���kԢ*c�%�,K;��	/��_̗���ٱ�B?�����@����0�Q�`��=�Bu����٧��V��W<f�lp}ny�x[���wa\�=9u����,�͒�q���N?kD���,�$���ό�;�8|c��	aᛴq�x�ȫ���Wt����U�e�`��x��@B'���
Ӥ�_H��^Gݬ,�B˥:ya��|u����[VNh��ڼ@��:�S��tq$����3�诌O��^|��)`�Wh9�RP��ϒ,�{�~Q���Wg�}S�����B߲������Tq�I*+h��c{�y|$��2r+y8'z�"����*��L�4��"�ۙ�E��Rm}v�4�K�k'��C���)r;�X�K�x�]�ڽAW�a�+��ƽ \d�L��d�k�^�=q�����k%���>��B���זi�(�}o8����EAf�6�Py���5{�	W�<?^4
d��������ׇ�����G�E����C�Ɨi�T�eqZr<���^�ŝ���v)/b����3As5^��"�!�� {��ura�d���bD,���_A�g1ψV��Y��	�g������y�R@W#�?Uq��%����O� =N+Ln���-��r�	���o���X0YN����Z�qq��hy��F2c���U	�1���Д��U��P�㝏c�Z�
W�L�ٰVm���x󚝞�'x`�����j�G�O[n�s�3SU�����W�שqt�ٯ�9j��xz�Z4�	r����lN���|I�:���5���.�"����DBէ���)9�O��X*���b�7������qt}�sHC�L�͙`;��9|2k)U:�t���y܎�Nq��ץ�@��@�7o�W|�x���L���Xx�_�\���Zo�G���nt,��J���G�QJ���"}p\	�gGO�,	�K\�f!�D
��� �V��ɲx�S���o�����{�[��k�)���*���+� qc�Z�0�+��<hO�c�/�G�q����W�����S�=[�w�G��v��D�͋'{0�2:B�n�[���#�=�P��'�0�P²�i0I�
J��C0�����鵯}�#�I�C�<?�F����w�i�l���:����i�r�]l���E�ù�Q%�b�.|O9��ߦ�� y&�dmf:���b�d��=6 ����`<n1JP�[V����YZE�#c����p�#�sŠGU���ˏ�BE��a�u����h5e�L�*�(�\��({��_E�v�z�=<��_�,�ߩ�H3FG,�����01�P�3�8����h6X3�+�%G n:4�����:���2��bOP��4�|I�
��t:�r"�V9)���(D�\��ةv������U�����ߘ��N��3ߑ��E��� A��#�t��v�� ���Ga;��)[������9�m}(N�8���j�S��W��;����f2y��(�[EE�K�����K65�d�ԾX����߼�s$�e��f.���˥����Z�,"�C2��s��eY��@?�K�
� +0�Z'�j9ss�6��V��t�/�~Y����h���F��b"v��2�97&��d�o�p��C���ӡ��X3��	�|�ة����ϧ�)x�[0��b-�^�>~��ļ{k��k�Dv�ރ���%S��Ҁ�wKi���g3/�^|[��V��|(�al2<����p�^c��y�`����
i�a6$SD|��Lq�m����G}c�)$AT���P�یT�b����_?Q�UC��pE?|�6��Hw����e�[�&��݂�I���6��~�  �݌���ǆ�%`w�2���hCG�VSL�S�oc�th-6u8���=�/����0��Hb`$yQ�CC�~�W��ڵ��Nk���/x{��}7!p�P�i�w��#�t�V� �� f^6�v΄qE��ڙ��zsF����Ý,��J��#'��ԈW�E �ݜ>�dȗt��<W!.�n�)_gX�(��B���dW�Yb�|���K%����z����e?�I�r\{�Um$����(�̞n �s��jy��"f���mT�'�Ji<�#���4ʖ�z5��*�^X38`Bi b*�-���"·���]��UC�ˬ9
��<��-�D0�y�R����or�3�I���
Q�ͩ&���1�"��؅�*����n�?U�2Z�"�w">�՛�{DM#�Uf��BRW�������9��4��R_s�*��L?�(�w̾-��8�JX�Ƨ�#��z�T�뀛PД�I�Yؼ�_HK�R"�GeZ"߰ �w�@ܥX'��r8��j)Ki�O�P���' �C��L&K����w��={̳@H!�%�5�m��o[ę� ѱ��,�l�ƨ��� �L��\7t�&�֣=/Ͷ7o�z�*A�I'�jLA���3���U�+����i���Ȅ���[|�����q�l"�t1qO�S^ X%L��t'͵�Q�)9�B�j�v4X�m\�� ���=h����- .p;�{[�+  ?呭��@g���H��g=ҍE��;=qA�6����#�>r#��:Bg8�~�[>��;ˣ�M	�3km����#Iߞ^��Y���JmiG�!�P�c ���=�8^�B��W>3�".S,Q>�y���ӵ{WϦ�V,"��2EFF���O�RJ:d���O�^y�6�Gn�&w&��di��X��N ����1[|`~�|�~`b��a-�eB�� ��p�	�Qo�':�'�L# f��ȂKa��`��7>�����^EL���xxi�޺KK���Z�}����k�+͍��gcv���/0Щ3�޽yU��SrV����OT�X�_0E�rr]�tKe蔛!���KT�c���ϗ�S��=.�c|�<���S4�ߍ��9��L�4���b����.(����E��|9T @��:���3p�q1 m1EE�l˥V��0Qp�������������K�_�˯m�LȐ+��.4&44��L�r}�͌kG�xI1�;���6�|Wr9Q������t�Z���6���l*���XO��-_��n����~1���ը޻+����E����4oܮ�a��o!����P�_�����d|�i���LS���r�8�Ը��+~��i�d~]bҔ�����ӧ���
b(�K9.����J1 \��F��_8?ar��]�O�P��(����}�0�X�� �:{*9t�#n��Řh~����==:�p����.�0� 4�>�*5a�_ےޏ��DSܹ?ҧ��c�g<������ivŽU��T�`��s��6
�t�72�<U�`w��%�Hs��ܽ�6j[L:���FCz�����V�A�
��XL�u���67tåRVo��N]e8��?�UT����Q��VT�^ȁ3�f|���(�EM�(yc��.U|\b��AT�W~���|�!��S� 3?.�N�h���#�z�M���?��%r��J�4�M~j��6�p=:��bdVlB����Qm� �E�w���Hx�o�ʞ��C��X�1�?[���+��/�Y
"���$�=?�#�E�3J6�f�J�X��ꓗ�U��
6�Эm��u�!���Xg��-�U�^����pw���h�φ�wh�k�P]�Н�wßWt;��&��Y����5c=#?`��V��ν J§�6�5�/�V�ӿR�_|�;A�A�� "%%]���F&AJM?� �:]����[�>��|E���H�;Ð*��Ť��e��U���5#A���o��ݔ����$��^������ j�@^�q���48g�F_�H_�`��g�=@�X�3��M|�����j��B���g�gZ���}�;�\d���-������
�r\�n��K��V����	mm�z#���aǬ��$S����{���^�@��s�[�PUd�t��D��N_1"��nA�ȸ�nэ�*�p��ՙ[AƯ�C�xx!���	K�/���$�:*����M�7��4�Sl\�W�ҿ3mo�&�>e�jX�&=�͕��ܜCT���+t�/��]�N/�P*���<�>�R�I�1�!�S����'�����-��a�h�߫�Lu�>���~�J�?A�'C�[�E@Z���Ȏ�Ϯ^�Dϸ��	Zl�f~���V��L4��� ����\u��'�h�E&$����E�䫍�oM��?�e���F�6�қ�{�Ҏ�����i��MH?w����}JY��W��B���I����n��7�0{Μ"{��~㎾o�]t�?�+��Iȕ����>��D��<W�$��	��A\\`�naAϸ���Oƣ�
[�� N]>x4�k.�J]��:?	jٵD((���2�[ݵ�B���v�`^�ՊbiôI镙���r�`N�R���������x����N�1Z�q_"6L�������5Z�F��f�v�ɵ��z]ѫ%6��]`){���IJ���03�{*����`�y��k�0b�p n�1B@D�";bd�����&Mj���ퟴ��)���w9y�F[2�Ƀ���`S�Fq��"�a~�����$CPBB���<p1=��oF)Ar̯H5� ���zvN;�(��s�����{��eN��z]�@��vv�*�ۇ����fj0�{�Q)r4��Uf�L��e>h����0B�(���	�۝!��8W�����]�~H\����U�����5�R+���ڂj��?Dq� 4��Sz��᫽�#�Ã�|�	��.K� �s�pW�iQ�K+Ťy� ��q�7�F �6I�w���p7S���n�-���#�B>e���ou�]]�j�L��_4W�������b0G�"��3|����Al-ܖo�zt����3�eֈ43\f��e���S!����[	�*���o���\�����{��`�n0�i^��|T<l�D4�%�G��om-���L?�����k���������޳ۜ�u���g�]�ϽPJN�)Wu7(��b"Ri��Yf�� ��(C��}LM�����.�'z$�`���hLF��dA��Ð���,�jG?V �F*�N�@���o0b&�iW��k��9?Z;w'���w���}�Fm]S���v!���/��}c����_`�˸|�2�fv��?g#nk�bҞ��I}�Of7_�q�� ���bs����C�����������8�Z\�t5Z`��:�E�~t�Z`��88��z�f�A��e>D]`"�ޑ�#maGu�U�o%����'),�c���K$��b��-�N�oYYS`�J%�όF%�e�0Ŏy���D��گN��wݘQ�J��)�����m�NM$��S����ԗ�C����TdM��B�d����%�1�2c%K�ױ*��L� "�0c�nB�i,��������}��1���{�s�y����y-�be�܇����`��eZ�.�qhz�C����h>��c��=�������a�9�3�c|����=[�ȋW��p�$��8{��b�6
Mr�K]�>>��7G�������_ܯ%�}qZ�HkW��2W��v%p\M��4�p;V��҆jbʆR�v敘�J�k�
%�}�@h�(V���l�K�kc.L����,�� L���Us�ҷB�	9zUd�~7�G��|I�`��"�MLRp5ֲIW� V��U	��d�p���"����:xِD�i�˦�J�|��,�$���=M��'h�.���e.����!<q�Y����֏��w�S�H���bPc`�֌{ 4bP}�r\�H�~y�;w��K���ㇺ��'x-G,�Q_|�i:z�� l��~�V����$��"�s[ ��!����nY�|�0w:$�q{S�;�y+'�𧨝�8�l���,'���/M:Y �/J�{�2�c2��sT/s�U
LU��8�dD�mw��V�T����Ɉ)�x"���Q���'ܡ�:x���kY�����Z�&귱8Z��|�K�Zw�L�P��V��rZF2����z"�e��
s���[���B�}n��Sw�'� ��	���=���{��W�WX��8�@�{�C;�q��z�U-�\3Ӟ��V��#�)j:[��G$�3]���*��-]�)�k�0�k�W�����|���ϯ�n�ؕ�~Ѿ�C�ΌZ�J+A��x%��ΰ���Fϊ=�E^��v<lb��4���1�2�J�Sz�A��ՁI_�#t��f�5��%����Dű��4��!�ϊ[��DA1��Ā��4��a�F�_6���]�wH���*�Q�::�z��3[E�Ep��O�Q��b:� �G�^r�OǭY1��Á��P����.�[��<C�/8��|Π*��V�M2���3�qz4=�f�iz��.�h�ކ�1�kd4��Zˇ�.����i9h�^�Its"�F�཯e�N(�`�!�R�z���f���p��S��T
e��ü�� ��@�K�>�%ϝ�vA#��c��Z#�l(��;M|��ӟ����m��䄿��8�z���.D��~n��.�����L��O7�]l#��L2o�8{D�n��+�����Gu7=����a"���A�S��ޒ3������k���t�,��!Y!>f���d�kn[+D%h�~<���yfx]�xB���Q��U-�)�M,\�]-װd��*Q����o�����]aw�^ybʗ�=����a1�<������be��i�Y�}����e��c���#�þ�!W�~�0�~>��".
�~��n�V>����}XQѰ�>��8��X/�#�ݵAoWf��Z�����[�mOCV�C�Z�z{�w� ⌂�O6��wkY��(p���A�S��7ɏnDK�5��)ϻ؊�����?�GqW�`*o����l�s�;.��d������ͅ��V�Ч9�ɜ��\�!���i��Q18��@[�x�/�KXg��ԛ��ֿ��]aL�>.1���n��տ�e5��t�׃�םdVï~����ՋBgބ�)M�[���藣CPgH�8�����`H����+`�[�Z`��p$�*�IF�97�ǖ�S̞��
�uD^�U6k5 ��/߫S������ą??/,+��M�kn_����[��|[`����l�)��7���WDC��ɘX`xX�k��y�;�]t<R0�u���]F�]F�	uVІ��h?m �N�ӵ����lT�0�n����"�+��HV0T�`�_@�=2�?�3{(��B�j�ՠ�H�n(�a]=G�ZZ�������q��_:��N^�&��Q�\g����F���l�Ĥ}�Go1�6�����}@���vc0.��(u��¨cv�jg��%��d��I�ɲv� �]��EQM��;&&��u<�k�zi ��ٹ��Y8�Z$
P|J����0�~A\��幼��3��Vv�,��<	_1V:�ֽ�;��%^��6����y�aH���ظ)@Ѿ�x$��l�\�"X>=��;F,�`����^�[э�ٯs(
^���3�N�#]����I�w��F����8d6���]w��'i(��~$���+-'��'L1E'̵�I�F�K��s��E��+
��KY�	���<��oY��Z�3Rj�
�l�W7�,���[)2F܆�bG���&&�x��������b�dL��:��^\x�K��{�;���|$��H��P���1pک�a����shd=p��Ͽٝ�d�$w]�`.Qk�%��+&y6��B�\e~`)~�`��Yw7��ܸ��*MϹX�ggk�^hO��"�ܬo��Jౝ�}J}���4��T(I��f�g�q&U�K�_��8C�~���m�ZXf��_���J������湃�����~����o��l�)͑�1����`Դ��K,q�:����Y�t�p�{�փ�xp��e+��`�ފ%���y�]����Ѐ��>�z	{��>`�����^T��Y{z�|��,�e!�+��-.��<�=z:�ӭ����R0.�}�$��X�(��	q��-?i������\��쩜�Ř���]�<O�P5��{��� 8h�r�,^_��%�$�ou|�X�"�=�[��on��"�)[��ߋ_Em��=s�肖+��6��� ��(C���f��/�k��7�
~�s�w�h�d YP���o"$�����(�үݪ���,Yg=��c�(Z���Ih%�j���`B�Q�` S4�T��o�p<"��Y�
1& ���"g�x�K��
����%��Le���i}��8��{Γ���ɭ����z�{��4�LW�OS�Hй��0<����_��"cW7R�
�C���e]ꀴ��#e�ڧi�_]��uUh(� �)ul}"�?D��o��-0�B�+>��s޾ބA�d��d�R�}7)uM�ؙ�6��
��0pJ�U������S'����~ ���`��ޛ�ߚŪ4K�o�3����S/�ie�E���{�[�~ȇ���hǁK�z���<��#;?O���/Z����<CU4�A%D��4`��__�S���(ʚ�����9�-��F�&af�����ĩ��� �T�_��s�<��}��P"Q��k���˸.��i��N����+B�8�7�eud�����5'�y�eW^��QSC�
I~Pf��܄ӎ��,V��O��e��.�n����}~$�|�!iS����!y@���qJ�EӃ��mo��I��%^���1b8�H.��8�"�n�=��E���Fl�_���Q�5�{;*~#S��O�p���%!Hk׽&K�׳��>� -�77A���Ԥ.�]��%C�؜L�hXE ���S�M%��+�hB̈́S�w&���T�MԜK��6+R�8��1�s�~�pl��9U����O��� ��^�cix�L	�3�8�@|�M�E�/���~ħe	GT��9A�S��[K��W��S?w�k���H4�T�lp{,y��A]���'�O�P�lmt>h.ӵ"���4�nm�1h��4Įq�Cn���CƆ���+�y!` T1\ z��,��Z`��8u�Kio�JÛ$�I��~�P�a��^t/���ڇ���\���$�s��@�������	U���H��T�;O`�� U��=��y�D��G�:;5��q��5��W�3X`�w��]m�m �5ܣ��FD(2��BI^.���Y ΅_�B
���fh����@�eXG�G����d`C ��C �#�<ݥ9*�
��w$��J��CY�eB��C��-LX�	���p��T9I'?dА��k�H���1����.�`.�f�dz�<�|�p	�&�K��SS��_�P��u��f��x�}NG�|�s�g�l6�T�	�
�;t��ٴ�����[��X��2�����UD����H�M���1܂�o�N��(�,��'��h���f�L��Jo��M~��C���'��#���2f
DRƛ�GZ��K}|S��k&D�o�� 鈍�O�m-� ��늗��H%�/�9?`Bp'��f��",�����k�JJ�2�. T��A��S�בK�c�GH��֍r�h��n��j�����:�(��/�
1��o��nY�?�p��aL�-��l0!��� c��G'��[R}n�&L�7����ՙ��˵5���4����N��F��F����D���
��K����n
hZ�-����Ҿ�;���'��(V�����	ᴴ$��·�0rYΥ���������xT=��`JK�s�6π	Ҩ����S�`y��U��~Ϯn803�=�Z#w:_���B?0Ŀ�����b�~��?ׯ'�|K�5��#q�Q��3φ�jV#�-�}�l�wc6�7=�Mp�.ڿ��U匿0��$���o�5�>����3�S=k��tH@-?�mV��>�(�aҍ�>E����ȅ��)��T)N���y̌<�s���k���s���[��3�W'O�̉�-��_-3��{�K� %��"�\��u�
�H�Y_�gk�!PV�/��h�tn�cТ� ��vq���E��?��k����� +֤��ȁy��2q�p��^w�<��+�l��ݿJ���E�=�Խ	��~@�N+�D����%PZ��qǩv�J<�
Y��K ���c��>	P#�)�E6
�7�e�����u.��8�Y�y�.�$5�/�c�c��&3�q__�����r���f+|�����	) �̻ �!yQ�P�uJ� :J��t�{��A����[ھ�uϋ%	ʘ2�薖�����[�
�e�/T�\�$�%=Y�(=f=�"Q�h��D���(�e�o��D��8~�E�0Y��B�B�� ����0\�v�*vW_��
��M�CO���e���d��8�C��1ϥk�Wh�b@�m����Ҥ��Q5���HqMѮ3��"����dl���L�lH[�0��{��>��+S�&H���4��������::סu��wy��B"��E��$�LO�{���\Y���`��Cv�ͅ�GJ�< :V�0�ϗ�J7>E���N�b'�}(J��7�+q��BϝvM�I�0�˦{8=Ε��gNe��n3V�70k�ZJ�v���E1���R��Mxͷ��u������፪��ͪC��S�&����i�i'������J��w#X���r]��Z����mj��(��[5C��F��,,���ě?��#��_x��G��ȣG�B��̗D���z �K��� m���2Y��w�Q>�1�Fd�����R������5��~+����ӰMK6+�3?>-v���VsՊ ����rU���(�y���3�O�g|5=��w���woc�]��)��D
S#w[���tMnő�n�ř��$�f��=�m�J%�b�ދ\���ߜ�ߺd�S�����0"�ؿ�D�)�������:~�{������{L*�
uZݐ�p�e��|�(�/�]��r�	Y�W��{���߀vYN�%i�J��^@/�	�C�VثĦN��d��z�_4g��&KG���lw�c� ��R�m��M�T�I�����)��{��A[�����7'�klZy�V1$�:Mhs�G�?���"��f�ы��Os��&p�
�$v�B�����#���������O4z�elL��yiҩ��h5IA�Ρy��=�I�K$������:�;�u��3e_Q�d!DS3k?�	.���t
YP�0�M���B�0:�"�fQ���=�M��W��Ʊm��Mui���A��S�K�3���A���o_0Ԕ����|�����/��f�	x�tP�w�ݢ[mB���v��
�o?�{��2.3xv������l���]���y庬g�ھ�����������S���+�b����
�p��Ý)�����-0~�1{6Y��w�))���
&����D@�����)#��0o���	�R�\%��W	���A�pš,�䖔�Cк�th4a�Z.�ў����,�f�w��վ�}G����G]U�U��p�+�|y�#<�<,H�w�`��9�����m0V�7��}�S�p���l`�T�l��)����H竲�֡������9vg���ּ�?n��U?����q  ^U��-�8m��O�(�b��^�t�p/g��I:T�s�2H��U� ���;NӖ��o/�aG�Y�W� �ќސ�}��[� eͿ�l���G��tĻ�Oak��s���"Z���4�f����՚��
����X��8����{(Q�^��/�k���b�s��P�Ҽ9^��
�R)��Ҫ��D#v��7�s����Ic���&@rl ��iW�:�X+���$Nh�Ŀ��F
�S%B����)��B�V��]d��᩶T�>em�AwA;�F7��ã�q�ѩng��H$����o%zQ��э�>
$+�;�U����lȑ���(t;��j-G�2&�}���7f�'�����<��L�����
J��9 [�^�*���'h͖a��xr[��-M�Fڄ>mE���%s
{��6~|[�����uIb�΅���aW���x�k�q>�?q��<���M�4��
ӧ_
X�+@Ó�l�gr~�t<�(�׸��S����\���t�J���:ݾ��V��������mĳ�9�K����$�8F_i��-i�����,ۿ��F��ΪD�|�9>ݬ�P�Rp[�
`� g�=&�E���W,P�d�+s���'x���S�L����
�?�a�)?Rf�����a���C�*��w��Jp�I���9�x��3�L�2��F�����	����`��Ru+� M����DixT>�����E^�׬�P�����}����ZM�z�K+MO_XS��_"o�+���O��a�Կ�~���6�0�jނ���`���W���o&��,E���ͅ
n���%X�` ��E�l�,��}�*�>��Mg3���3M�i�J\y�W��&�7�F� �%q1F��?����@ӹ��&�	��qnqᔌ���Ǖ]�w$lU/���-f��(���no��H�w�K���cgsD�T�\�(a8-���c��V~����]Zj��E�`�n3��tQ���ᣏ��p�'S.��E�댛��.V�^���v�\�F��������u��*L��M�gf#G �#x����xו�)�}�:�N��������2+c?l�ε��U��;]K6ʮ7��)���~�L"x&_��HR��3���/Z���7�]�����%�}R��[9O��K����TV�w��7�������䧟A��J���p����������2fI/�Ѫjɺt$6�ʽ�a!�| nj��xҼ�ڃP������/ c��P��g
\��,��J�|�5w���t�bo����*���q����:�Ѩ��H�D�U�.�6_�vJ��-��ə�L����۫��̾�񔵏�s��n���Oeq�Ϛh,�N(��ܜ��s[n4��gΚ�����E\T��fR��፿���>]�f���g�|��h����^1r�9 6kr�h*����Ԁ_;��9#�Z�+��eMM�rSEwi�0�������2Ȗe����̍�`�%�;��°n��p m����6�~�7�.���݋�Z��y�EU�h�z2�0�tp����ܷ�˄�l����d�XO:�G �G`l�Ds��YM�N����mV����fAH}���q�?-kx6:ӳ$��w�qg%R�sO�Ω�JX&i^v➸�Y�U�������d�?,G{��oX.F��g|��K{j�fFq�=��G�v��p	.���|a�����S�߿Ij*9e\9�v�_�6ω��|x�]�䂒}���ЪDЗ<0�e�����U��9!���I�r� xF�TT�?�]k׉V������L��aVLw��#��L���	-�cc��0�]�o�²���Я�R�o�<&B�Y��_��u���h'W��~��*�<�=�KBy]:��bEɭ/q5
tp��@^3SB��U�,<Y��a�/-�74h�z��҃{y�U I�6�e��iX���#W��F���e��������Дjf���4�W�={{�e���F�\y�������l��6ܵ�+Z�w;�KH�}~K ��tvMYP���o.Y���E���l��;j�'K�쥛�A/?��@77�ş��E���G�u�g$b�fѦ6��}����v2:͜����#�G��T��;��#k�_(�X�y~�!��=g�z�z@�4塀�U~�β1(�bɭ]Z��n��c���PS��$��wv5�-�`�٨k��K<x�(����V���d�Ѧ�4rb��'צ��N�=�<	���Y�V���P���m���o{ ����k ���c��t�qͭ���m%���W9b�?x7����q� ��h ��3#��˲�w��S`*�e])��*7�33O���[�| S �m/�|P�tT�{�0�_�$�?�����5>*y���
g�Պe-g����.{	�p�;BO���P�oXR*�lt�Y�XhT&��}�[�����|�Oޡ�y�"�h�J�*�E���T�u���"ZU�Y������G���Є�~�g�1��{�Јxs!>T�C���~ܴ@�8}�}I��X�!+X+~�����As�� �ڔ�������u��bG�S�ޒ����P�F����Vcje�#Z]���C���k����ǡCA�Ņ�Td��0 /1�Aڠ}�u�o2�����GK�2��ׇM���T�j�G��f���P�)O�x;�?:G������6GA(Vb�X��-��v|��`�+�/��Ε�d�,T�����?<�9�L+x��Wdؖ�/��o>\���:D��F�1����?'Ev]#�m�	}#�ܜ����x�V�yz[�|`�^ ����b�������E�ߜ� �BVg��i� �^�+KD���f���O�s�ٷw��J|E�ڰd=O�t־��W����Eqϻc�f�_a*{6Y�Z�'cK��ӏ�Lu~�6��#?���"�������x48J������#x�٫�Ԩ;etT���^T�BA�	�����ME$�f�5�QPN�,w�^��P��C�D��u%��-��v���p=��T1����r��(�}$�r9���D��W�K�'H������?��(t���p:�1��6��@�F��t���ޛ �5AK*�-��1a~~��>���V�m�Is���?�߷[]a�Wf��Yv�{�
�Z�`��������U}��p�gYc��*Ӭ�	&Mq�I�4.����tTL�A����ff��"�j�XN0�y�?��l�����#��������oG�8���睒l">�6{���{��������J��fb�\��o�w�z$��	Y��z���M�j5ƿQ�oFxQPR��ҒH��~�[{�����m���cL0(,�����
{8Kb�U�ݲۼn��i���I\ƶ�y���:\.����]AG�~E�� �/�6^ꢾ7�jI\��xr�w��k ����\%MKG�υY��$�82�Q{+tNZ?+3]#b\j�>g��{�3`��~W4�����~�2ʾ]�~������������Q`�H��I�`���Ek,�ݾ��I=x���X���~a�6�E�F�ky[a�[��+&�E+���� �_�81&
����v�h�DcD��>�B�v=�+w��DJ��ӻU����W��b����d�,�������Cd�T�	�D��g�FPL�wM���&Lez��.i-A�:]�̻��!$b��|Ii�{���鬗X����q7G�����<�gN��b����~�=���S��V��s���֎�z~����`&���'��T��?�p�� 7 U�o�u����/-�VY�4	�|f8>���Ѕl��m��QZ�X�]��ٯ^j�Vp����`1ZF�N7$�3-�;��r��f��W�'���������σ��� �V=��$��pu9A�L0�Xۇ���:.�x����)�N�z�I\+���ݯ�����c���[c�EQY᥮���wA����pQ�.�2���_��D���O=bɐ Rc�Z��,�h����z��Ň���SӀw
�UM̳�,���x��_���b�7���#�ʬ���A���~*Ǽ:�ĝ}�`��)}�k� 2)������x��l4k-a} ���H%��� �����8#܎�����>4�%�N�y�� �,#ګD���X�W���F����~>�`����瘧������݁ ��XMV3`&�
e���KKHH|�ic�~�yN��x�1]*�Xp�(�c�%�۳���X��V��!T[�l������8Sш+��W������G �-�I҇eχ���m�yC�#�J�\��L9����}F��AN���X4��E�&�Q�R�hy�K�ܖ��ڥ��t*�;.��� kM�>��(`س��ϾZ���|��}A�0t�~!��=
�>v�Q���I�"=�9�n��j�5��P���A�~{�2i�����תz�m�� �}��"���>>����Z��mhx���E���r��)P�/$�r���!��ˇ�����lh@����L�֫f���Z�Fs�� �8���l����j����f>�PO����W_#B Q�U8��k�\u[�jxQ��vc�_�T؂?���I�[]@����Xb������bx�?F�G��T���B'����U$��(\O�9b��j�
=%��������blb�%P��eF��}��"�$�5+��'��5I�yM?|�x�3Q�&(��=�w�I�ʻ�2'e-��*�>/����P7�8+u���7,唦���Oc��t���g�c9ki���g���['ɢډ�xs�	;2R4xO.Wy�>�)�)[��$���YwH8+�=��G�;�OhCS֨�Js�5���k�Z�S�e��}5��bn�r�Q�3?��m�N�c'���,�4��M�Dt����&�D?��i�-NͅF��� �Ō4 n�AM-���G{Y/����<��+j��P��pq�ޅ�Qn��d�t��YR��?�R�+�}�-���8&�T��]r+��]0Wx����Ǔэ^ح"x�"�oQ/�oو+wc��_�'���~Pl����2K����@��ؙ��f�T�q��[���w�G��y=%�����p���_*r��N�0lSln}t���nqc�v�^8I;h�&hp�80���v�h㍿5a^3�-{����^z��� RN�'3��L�DD�����WPj^���u�R˽{#I�^RG~�_;bV.�.OU�;*N�1ؠ�	�����D!o+{��|���IzZ&g�9�v
t\a���R��/p®0.�7�u{���sn"6-�����x�x��X�~2��S&���7�X�X�	�t���M]T���;���Д��t�����#����ٖ�v�&���F�κ�`�{J���(�pV�p�v��"yƃ�����-D����`:Ë��q���W��e� i�Ep����e���ʱZ���������0Ԉ�,L��!�1���h���uMA8��}�-�i/�Sd��$��̌`��k�ޮ�v�"&�g"���GHƯ�{-uU�CsO�}4\�ζO[{	�(E��z���Ѿ���G��(
��7���]�e��zX��~4#z>hCu�v��FLK�K����R�^��H���e�k�7�<nz�Z�"�IՆ�9���_��N��_���D8�~?�"�z,0���h)��^_��YI�����g��07LQFR�(�D;���8 )�4q�y�t�w��QyA z�C|CQ�=˞͡i���v&^?�x����˸��?�t˽B�v��ƾp5�t�px0C��qp����]$\�W�����o�V������YډX��k�V�Zf�����o��<�l�Ѕf�Wi�O�
��BNPaBp�Pi������m��$���Y���l�-�c���6^gji�`Ƭy7~=�N�$�+d1~���O��A�.Zr%v�N��9����o��Ú]���_���	c)���LYd�=\B���U��)٧ɢĦM<t���p���y.�%�;����'�Xt:J��`0��Z�k��x͌��H$5fB�B��]���s��w�455-!9���{����:6�_������|x��ޮ� q��O6�� <���P���,w\³�Is��m&�ol�W�'z����-���o�ܻ���;l�9φ #@�U�#:���_����_���B�ѭ����	c(<����{���耠1�Y��ӧ�:������l�����)��ls$�t���wo��q�Z^^~�?F(r�{���@$�<�'�r��j�^+�~�]:�논(ç|Nn���n��������Ǚs	��P+ �C��i�p��qn��+�r�=�+I{2���%�f�`�­�-1��_��#�kbN���Z��+ˣ�	��5��G��;��/G�&Ђ}Ч3,m�-t9�����=�Z�d��h�u��\�8}[0��8<P�B.m3G�3��5L'����- ����p53��V�UW�b�K�6�����
4��F����.7 �Tml�*>j�}��ZY�z� �r�F{W]�t��әѝn��_��|����÷�}ss�$�<}�o�ZG�?5ީ��/i�R0�5���"A���QPL�?\ָ!x4/�ΰ�S?NN���3���4�6�@��޷C��E���Z�*C��k��a���V~�vY�L�ӿ�ps-���:`�B��� ��oHs0�˼�Z���/�w={kY����d*���`���]R��2*�V�>A>�ݠ��͗7�l!@�R���K�$"����k^�u�K 3M�@9����0H�~>#��������g�����i������}����	�</�7����J�7�'w��_�CK�^nϤ%<�����������A	��?֘,��,QVkP�Y$��=�ϓ��������ߘ-�����/�< <�z\�����&�Z�m�Vw�o�k�D�aK@D2�?Y.�k�M�W�;�;�ѬǛZ�Ѵ��@�Ԥ���B�Ⰽ4���L\�J�"��㡲�.؟��b�d��8R�������e'��vsx���G5ͥA]���gG�����P�cx�})�u~��U��<��#C��_^c�<�_T���+8�.;*�����rKe荎y�G=��~"�{�Q���H.v<�"�0M�H��-L���d$k���X�9�i�[��O4�ج'����٪�˱�:E�.v�]�o�
�d[\X�^�����U�ƃ9޿s��%jhL^���E�U�t|��2�\-�Ju
R�E�9dcrr��"?�	�<ſ �R�2Q�LM�z��6Y(�׎�D�)@�AoO%S$Y.W� Fu[�bK�b��+�Q���@Cu��y�goo�ȇ=c�YZ���̲�J
�з'���)��M���W�I7"'��<<��*t9EN��������Nت�
���(�4�1v���WW��)¥~��RPK�Rk�I֧뙝��(z�����4�C�5$h'ީ����@�ߧ`b�+LKG=M�ߪ���V�'(�w7��܀�}P���Q��%e�D��I��6�C��h�|��4W��.�,�1)�V@�p���zԒs�z��(&�M3Q�i��	^PPp��h�i���(��l9Zƙ !��"�.�w����)����;.5O�y�6y��������L�h�qg��7�ϻ���?��_X�k[k�َj۟{y;�B�C��H:B�t$$+��Y�#^����d�{G'�d@@�� hB�h�\\,�Z�V�?s�ȴ�B�Ј<֍�0��i$�>P[�r���ϐR� F#2�d�u]
&֭r��"6�k(G2(<�:�2����R��[^j��?�q*��z�}Q2�F�¶RΖ�l�m�rU�g��Δ�s@|��i�$C2��/?'���˼}|��V��?�x@P��}>��H�M�
�%����Y%ۦ�$l`�L[ĔN��j�o�~�GGz��o1���%���>m�C都�r�q��E\�T��"�/ߢ�?[�Z^K������/�A@��W�*u��6�֝z���F�W�/H�j���l -����0��������v��4�^/�*s��Р�RΌ�(l7��u��R�@�E*�R�#CD5|ɶR���H~�ZZ-���ԉˤ瞞'�2Fs��+M�5b���ϖV�R��P<Z)j5��7���j'g��/1J�#�����9���Z��Ѹ���F����y��hU�|�|7�"DA�M~t>
|�1!$���}����-�HeM��&fVt��#�y|&�u�
~.����&턪#�L;Q$?��$�$��u�饅���u��!h��S�f_1�y�z�8d����h�<}{#E���|�8���:Pn	�0�1x�K�E�=o�۸�{l��Z�GH���U�\!�T��Qa<XI����)+:OZ�`�@�<ws���/&k�sOm���ᕴ~����
{Gb�Abuaaa�r�
���JJ)kGc�CX�Ud�LI0�˟���A��v�c{����'����ܡ�}�����(ǀ���kpr������ynr,dl�k1J�*
�()F�X���ʜ)k�㏘�O�4sof{֣�*۾�D�}��ѵ՟	����|�SR,��p��6𛐃�Xh�5f"t­@�#Q���q�	�O
�j�S(%3�ލ��W�����'(��.yyJX7�M�zl��}���ߟ���o�� X�`�Bι����Ec��LPJ���Z
T����*���K��e��򦮹z�m|�lo"Q`Bz�s�K��n�F*�|�)��G�h��
��:~r�E˲I�?�\[�ޏ���<��Pj����#b�7����~/�r�i���K�NW�_r�C$��]k3�C�H?������0�m�����m><h�L�nU��67C�	'�BRO�\j-U^�9��({^f׼��pт���y�VO�5m�D꒑��[j0š�m��t�2Q��` ��@��&2d>ڀ]m���������O�h؊��E�Yl� �p��),�޹)�j@GW��9*C��ۂ�'<�5]pÉX�w������JGX��v��@]��$���p�;1ĲM\����� M_�F��g��w3NW��Ʒb�'��DQ��70@���D�Q�T�c��^��ݜ�
a{��q�
8����i�c��E���ⱒ�xS�����`"�k�M�����^��P��JM�K�T��@�]S,�ۛ���1A2�O�>�5O�i�?{��>}%�^�����.7���Yzۈ<�z͒�=���*t��us� �!�R2tF�X1h��(ʖz~c���b�ﲟh����#0�G���Keü��f)U�$>�(��ve��s]���_�覩��B�6�.��:�LQ�y�p2+)����4���PYn㈴�D�8���W�1�+L7<��\���b���grAVz�#�z�(��9��Jx�PVIv=n3�f�*Lr������ىEB*)�n���.�4���MSOg�	C���8IbV���e�����OV~R��{��Z6X��B��l�I�f~Z�f���oR��(:����O�ڱ�q����#<�]F�e�i+@,vTl�.��a*M*�M� >��!���hE���P�D,�b�j�lC�������Xy�Z�yK��HB������� �ˁx�!b�R���VbX#�����I�����ݪBg����}pl�&ܚ:ߋ.�)��Dx߿wk*��R3qKvC�E���l��&�TH��ohC��p��:��2�xr�ro1�f��qT���)�����<2�b;6�/w�v���ݯ}*ʝ�]|�b��bƯ�H4�s�Z��w�p��ynq���o[J�jiO��~kZz�eF�w�*���	�_6 {Q"HIv����0��i��?|xFލ�Nd
�h��$�73q���]wÄ�0V@>��MDE&}��M��(*��0>5u����xM�P�i�~��n-� ��zk	9��Nu<�{2�^��wm�qzz۰�9*F�z�����x��V����y�7*U�v�
�<��-�O�e��[d2��$^�K�	?]��>M�U
|R�Ym���P�F觃E���8堑�\��3�)�l��<q1�ʙ�W�A3���m �}7���o��w]����6�N��Ð+/�Ȓ�	���dƖ���Ig$�0�"��V��Fw�O3��B��9�^T?c�WX(�"`&�t@Է0��At�P�����?$���ZK��cU2
��HI��)ҫ�6pޯ��D��r�|	ha�;�{�o���$I���h�\�פ��?%���<97��M�9IÕƆ��er�o������[&�>�j"���n�j�\��Yx��_8��5�)�w�١(������X3wGT���S__gB��ɮ�.�jT�ج@���ܨ��H^��3w�[�ʇ7�����y[Q�h����O ��]�;�-AC[B�1d��Mv�ϸQ���������I��}�s91����4�f{ʞ�h]@���N�f�÷N����_�5y�Z�����q�b�+�_�L��I6�߶Ec�BkF�4��沶����)��X��Q��i�/@��{��V���Q�����3����Q��_aj��e�&�L�WaI��3p�϶$���'������T}�X	�F��wA�nC����XK,|��,(X�e�倇��iî{�Ⱥh-ˮ��dS@�C��+�4����Fo�(�(Ռ9�J=,l�5�|��,�ٲd�o��{�� 0�X�}��}���rbO�k�����|(#tS�;3��Kp���#�]%���n:<�����盈MV�V�Z�!焵뵀�%PJc	�$h030���V�����n /n��^q\�pe�*��:��`6k��m6�%L@?�O��e5@H҂BҰ�U��iPt;��^�wF��8�����F����mW��u��N��!j	�������@@\G�(��d�WȐ,�42�j����'O��D��Pu�>�te�\�$��Du�)�n����5��2���-`=,�7�|o������OA�����X��[oe���֍
Q*����Da�Ice1�d�4*-
7�mH�(Y��diȒbl�d$�i,Y��Be��\�}���<�\5�\��Y�y��y����xǷ��|f�2����*>]�����IE��8��֧����!�~��&I��H��1�=jY2M��Y}b_l�s/Xj��H/T����f��� >���`�3����T��Ћ��9�/9�x:�dm���=�_�b91���6to
 `���_6�G�ڮ$���������=*�fF��&��1Ļ�o�������jd�!��j?b\Ҫ��l N���DX�J�����3
�I�K��Z(C�N���R�e%v�ƢnF����?#ث$/Q?�Q1�ԥΑm���쁟|\�z�Vj9;~<X�>�MA�Y�������d��������Z4<����
�DN����d�0nR,ξY�Q.��z#@�_;�%�Y�e'�����b��T�\��)�n�u��.�Xk���ICDv�k�/���7������w�]���`A�s�uww緙p��v[s7����	��g�F2St��Z}<h�z�a5�����d�'� ��9��}�v[gk?��i"J�͈r��+.�s�0�^<��$0`�~���b)�
.ܸ��������E�}�U2�A3���+t#8�o?���
�T0�E�)ݤj��r��v����������a$�p��]M�˕�5�)>������cL�g�)=��N kS4����A1��E����>����{c�%c6i�exX
@h�ԓ��RP�}ю�b���uu���;���TK���y�^��0z?Vp;������־|v����H턉2���W���^\�~�g!�����/ˑ��5X�ղ�D-'C��	��#�� �H�©�~6W���N�^�_�z�f��b �,C��W�ش#$}��*B9��?-�bп&A;���/N�9��۷����Z,���Q�s/�\���w2���<-�E u��t�g�P�<���u��2/�B5��ݪ�O��@�G�vrEm^U�rvUO����
��nl��r�ǥ����fB������}�c�D����Ϳ��f�:������Y�T�%+5���������4#�'o��1:R1~���ˡ^b��М�߹;�1����_�侥�p�>�U��2ٖ0��Y)������(?ϙbG�_���
w�l�8�!��(���e�!8G}�p8���u��>0��m�T�k��O��X!�o}7%��n��h���W��N���p�(�Fͯ���xq|5آTmz�C�Y+Df�N���9��L�5�?�AG�T�9������~��+��gӟ+�L����S��^�1��5j�����!@�7�1�d��L�rY6F4��ty���a��U1ܷ;{�Z w��9�Ӣ�ճ�
�_E�$�����1�K]���5H-�<h�c!�d��D�<��_����3߀rg�L�a"��3ߙ�Ge�|NЀ?�\���f�d��Tda��!л�D��2��Z�� ��೉6���^˜e!�-^�8j���?��|�0�NTGZ�y�n˨��`�Ebg�鏜���l֑E�L�%���1��W��K���݀ii�H���MV��u��6��>��u�X8
}E�q']ȼ&\i�'��b��n޼�����h�Z�O�ɰ&�Q�h �]A.�+��
<���S�d�G�r��5Cs;�D�����*C��i@ %�n�d��C��/}��e�u5�@]�	�m	g(C�,�+j>m���0�
�tI����F�t�>�p���>�渝]���5�����B==JM�t-Q�\���TM�7�ꋌ:����QS���W�\�Z��y�s�w�R��m5��+���
%�;F1U�o[lr�pQ���g�=S���/ux�E��� <��xX������y*%�Jx>����q�okY�4L�+U���^z$���dϭ��=�u:��Y���2,���KR�gTft�W��Q�1��{���9�:js*#�ܷ�@9���q��Ly��|����Ľ<��eW�X������wl��R��F�j�a���~��MM~�+��Ļ���¢φ�������*tPNo��?;_#Ѫ����j���	�@S�aK��.+� )������-��vA���zք�~U����E	?��nf'��l�h�mr�LɆ��J�g,U�`��s�l� �y���W^=�g��o����F���6fę��>��S4�u>����+κ�h���)��ۊ�zм����tO.g&�`��R�P*V)��Mv/�-����9�.�0���D��<� �l"��%e6N@�4�$������Ԯ!J��Ĕ� �f��>ê5�6#����Qr�]�	��CM~o��<m�3�6�;A��*u����ӚXeM�A~��|���[�{�x�/��L.J&�l���h�]�,Ң�Z[E0[�.���o���=�E���bN�bd�;a)���zw�;|U��z���Hi�^��H(mEA�&;�;ʀ���0�~6nnQ��+���ej�x͵���r��Ȭ���ǢE���8��ռ)A�R�vmdm����j�Xx[$:!]ȳ,��E�s��AY8I.[Z�<�Nkf�e8SA�	k~�F�S�p)XaRᚡzC�}!!�rUs�����E�����K%���\Ů�.��Aj8#����9%q[dy"�&�+?:n�w�F騳��� B�Ą����.�d���*'���KtS�&�q!(�i���V���u�� 11s�:G���ƥ�/Q=8Or欁�M�Z�CW��P�UමF��c̥p'_�'��;/μ�鼋
�Qԩ�t�{be���u�tF���:�Ih��Fo�2�V_S��d��fff�w.&�=�b�z�J�*U�L�@K�Ǣ��g]���6�n�gW$�&=�f�&����O 4C8�q��[��9��`�a*��E��Ig&fpR/�TA�0��Q!��|GV��bڵ�A4T�zPk�`Q��轃|�� �7V=��.y��X�0�3,����{VVVj����i���N���5D���%��̸�qd$v߫/���o�ƭ�/�_�|����M��V%nL�Wrw������o�Z��'�G�#��j_|�|[6�v��4�_�t�<�$��2�\閟��c�K�[�i\����xu@$tu�̎4y|�I�q�@��#�L�3��B��1-�x��B��-������hE�jӼ��nɎ�.D��2�t��B���J�t��� C�ވs9K!�%D��j�t=Cڦ���T.�iV�'���n�vX�b��
Ѽ���p\+����O����hD��]�/�l�|��ؓ�y���D.k`CC�_xX��
F��ݲeބ����
!Sn������J�g9C$:RRR���69!�խz�Ǐ!+��v�#Tۃ��~�P~ۘ���X�r�.��m���ZW*��bcc�i]�5�w��'2��{a��`Ժ�i��������^q?�i'}�{���Cgc	�GD�� �~r��������%6��<�E4e�'ͯ�X^�83_uR;!Өtǲ��n}o�G��΂Ϻߪ��Ʃ�I�Q�tuu�"ˊM����h���w��}O��݉
�/��g'c�S�;��:r���$�\o3��i���IӃkb
�q]�[�銬?��}�T?-;�z��;M�����FFd�QO}�e��Ev�nH��w�wҁo�~~������ȵ�00�n53�9������j���������0�����b���K~�?�#=�?s�|?�)�aL1�aO��,�|g�MN�k�]dW�Rc u���[4��WH�Y+�J�[��TL��;X��쫭5���{a�Wm�։�Ýu�o(&dJV:�]�
{@����R�A�����R�Kd�Y�O����7�Jb ��J�96W����r�%�Ҙ�wyя~p��MU|B�\���Ѥ5���;K��",)^��}�� 7|f���<ް��a;XD��U�{���UdOJ3��.��^`�i����0TY'A1��.׆��U��+��6 �y����>�5��?1��Z=�0�}x�s�r]�������H]�R�6��Yp19O΃��$>�*��g!���PU	�ת�j|T�"f��&�|��Љ8]+��Z5�'��3�z�v����xH�2#�5�O���CL[D�E���~d}�XmLP��*}DJJ|k(����՜���?�	�j{:�t�֠���A�%j��W��ww?��h�������~�y�3��͛��M��K�ن]v��c%��'����\U}�����`�M7D�]��f"�˼�݇��d5�8�`�%[��i�ʞ����G�r�J �����d��,X<W�ݓ�:�X�(Y=�6r�˧.�'1?q8�Xy�*��>����i�Vw�]o��H��Z?;�S=�KMn%6��-R�>|��#�����1�h��w������n��YY p����0����S��d�b(��~$����ض'���iK�E}[Ԭ��aG]��p��s����;�d9 S�F�h ��l!2��5�&wO� ���yc��y��#W���,V���@N�R��(���5�/X5I�}��uk\�n��S�a��Υ�I$��pw�O�E3�ZY"�us�Ɏ]��*���Y����,���!�m Db���^�ٓSe׮�70cZ���3�Y��j��HϚ�`)p �3td	j���:BԚa�z�_10�q������I����[^���}�(lhG��dpz������ �T Xp׾9$t�Q^�%|BE��	��vC$|�BB��\�\.���4���G�KS���D	:uE��_8ܳR�z�ﾗha�����ܟ��_�����F\m�m�^�~{\N�Y&5n�������x����d��技�����'}���Y]����=A�7�?~��p/�p<����ي� �XT���b5�����Q��U"o?��W��=6v�}3�'"���u��vҎ:�^,���e�#3��6�@�_�4Ϥ��#���v��	��D�!^��ߏ�#�2s(������^�l���6���E�`��Z�F���~bApҊJ���B�:���0˭<\����
+�	S��f__2�L�G��Եi8B�~<��j(�a��ۍ���
t	�A�t������Ql�?���;��T�(�~����ϟ�E<77�:�]=׫�Ϳ#"�;㳳ď6�O[���ٹE����$�Aa�s"ͥw��4S�������K�Au�l�>�w�r�^ˈ�n�a�
W�&ϡ�qv���h�%��C o���T�ͽ�#S��7}U�w���%��9Lk{NE@�IH�J�s������v`S沊��V��mu�[��[Ws�'�'q��b����lVū��'3Rd�|�v�oو�9�sʊS�Sbr}��փ� �./	ˍ}��w���$��@����+�[�`�����0wR�U����u/� �9ߊ�����]{rp$T
�=��?���<w���(�W����ll�@O�bу����V�6j�
	���P��uW�r�������j��ٛi����:�5���v03e<I��雿����9�:����r�TJ�O"p�k[����X�MN�}�V��>�T9�a��`�|g�e3g��%�=J(��������n-�&=��1���Y�:3ik;�XX�'��ɿTr��u�;��ם�3���ؤn�JG�ո���������k��.k=�-�M
m�%�m����<'ƶI������!�����z��w]��hڷ��m*���h��Ρ����w<!�~�e:}��UL}5|_�Q~�1M�.�f�-z��N�c�-�HZ�X(�m�u�lq�����o�W�%�_h�O�}� 	���܅5!x��">`�쥋G�օ�5X4{8B�jɾ^�����.��Y�G��KO����̝��4����:3 ���Z�t�M�B|"��t��~�v]�Q'�Z����mb�9��+����)��Ĩ����O<`��ї��ېQ������`�HT�7��1����V�J�Isr�7߀��׍NA=l�58�ۖ�E�k�\J�M����i� �c�%Yדf	���$~��-�K���^a�f����i���}��faJ��?<R2��x"��T�ڞ�G{5�ܨ���hf�r�W\p�iK7� �*��`���y�������6�F����u��'��;� k��Y��D��QP�F��mZ�K�LReW�0��iaϽO��)�9���ā�Z�����>a�Z81�v�=���x�6�! �ɲ�`F�rRE��IN%��7�SI_qUٞ���W���2��1�5���ju���+* :���-��g!�q���.A��A���f6I[����<ͯ��U�ְ���_-����z]��s=̬Ad7՟��,�J�����\ �W`��ҷ,�.��bO����v=�Ή!��fg����v1V�a��<���E ���k]T7>혧m�����L|�e+�%��	��	���6��2b������< 54���a!H�ǡ���q�l[i��-�zD[�ٝ�eEF�K�NE�ms����8[�VO �ec	����T���\��ġ�tn_e}���g|�G����$��ɫ`"����(�Vi��TD��)��x�i<O2��w�}�QŹ�9��h� x~m8;M��{�Իi�0�W�x��=���sY�p-����!V�9S-�\��d=��WKڱ�7Fbկ����ڛV�~;Y�q��|�T��o{���*����7��W�\��iU�x}svdS�������m9��𨩼��	^%������y趻�
���*R�&h<!��z��i4���.�qݖ�X��i�����
��	B��� s��*-�,�0C�	-GJ��Igj�AC�O_<I��r�칺�i�/T1}���ȱ-�MX>W�~7���	���4+�B== (�`Y��������i~��a�6�ϟ�;��4~��v������MO21�������ȠJ�g�n��c��7�藏��X����hbgN��l�$;�����7�f@���c7�lI�_{��&Z�}�dp���M�gm�I���s��x���;>f�f��ʏ�3�p�>�zqn����^N��h��B����ل����܄-+Q� �^���9b�
1s�np!e�6�|&mϚCQ� HK�V���H�-�=v�ǯ��2՞=��әݟpjmo�Ƈ�����p�/j��&gf���C����-R�ƴI��;���砱��VX<R0�v����sFh+�OzÖI%ļ�v��l����L#�?M	�
�6������w#���S������]���^�f���\�"HJ��/�0)3��J���dEQmX���GD�KO<*�up/�#���<�`W���AL�������N�"�NA����Bk�O�,�YO������E��J�~��ȿ̰A�\�G�YR�v�U|�E�5��@ n_��9Qבff�k�8����{z��q���{��5w4,�R���ܟ�J���6т�M�����^E���
� 5$��|��Ϟ"gw�4�Z�pn��-�;B
�-I);���&�d���-3�d��j�kof��S,u��b/F��i�0�H�����V��,�������]]��������<>����)u�^Z�K�f��b�F�����s.��7���/���5�6�����>O�c,�MQ��쳼S�9�Bd"9M+����C"��X8zR�",�:�$UK*�as3g�ʰ]��D�s�,9&�	��8��2�v�����I��CN�]D���>��P�7�)��r�\"��ֵkX��Nsj�U�6�Y�pk5S����－�	�<�&��2�dl��qWߙB�Ak����$/�Гc]�:���Y��5M`�	�2�*e��y�X�:㬝y��d�r��Xi$�e�T�@���_���+E�#��p�S�B
a�<�&��vpM�h�8�!�^*j��M��r���`��*NV3N��̲<�oayX����*�>E`Fې�#���`��Y&��3<߂M<�H�)h��x�<���'�j�����Pe!����n�my*"�b�CpB��'���$(�M�E�����0��"�ݣT)�&���n��T~�1KȽ�����93�Imma��p�c�&�+�!�"i "���=n��|�%�2\!rI��n�\X�aaG�8Y+����CĊH3QRS�(���96b�p��K{��j��U���Zh'�Z6F����qR	6q�<u�2�.v3��2�3�����#�b��8�°i�.�i�5P�Ip��ǛD�X�]|��v��(�B@ɫ�F���4�P z��j�7��L<&�F�Tf�J�9�T[3HZ5�7�"�-�!���t����T�P�b4�xju|܇���4�e��(��e~�!�X=�����~ON��I7f1H��"Ե6��y*����^���h��/�{�qRX=�i�x+=&�p�!�.+'y��&	���\f�/��`
�a}��� \�rח���E�����*���r����(�Q��l��"b�+J	��9_U�o#J+T݊�E��744��ʂ�?��qNyn�D�t�^�a)���
��庸��c�utthdY;>�MW遥B��ٮ�����g� ���Qu�5�*��k�ŋ�q�fl���Ί�齜�S������������g�G��'}U$T�v��]�F���h�����D�^���G\��T\�Ȼjg�I�ѭ^�CW`-�Ǐߎ�[)�M�0�;�q�SEp�3�����tX9M�w\�=4���2K�>����l;����T�J=gx�[��k�����_���)Ƭ6��pC7�6=��_d��*K��ʍ�E�9�Toc����o�o��u�N������������¼Ԫ��FIR{>��V���=�f�6�;j
w���`��Yҁ�Q�o�7f�0�F-Ɯ��Z:�<B�N�3�wkf�i#M��uw4;�NOF
	�:��(�(119e�z7�T���『s֓e�3[�TK�f����C�o~
Ж���޲(M�a@� �k:�ӟ�m���a0��۝�����sѿ�4���YY]�W^/�Mk}�����-��������ޏܛ�nW��ݹZ^3yr��GaA~����F �����>�W����Z��z�TO�3H�,��*�Q7��h�ŲVd3	$��Z��ӊL�I��>$x����r���Fy7\h;��z	ug�/rl7���5��]GiC��`U�W�x�m������c�=b~>^&`5؀;\�ɢ��W7ea.�Y�	����]�#���[�����9HZ$
�(%������ADVk___�T�u-�w.�0�j�w�,�Y�����/6V�lŗS��k�β�f~��d�$p��d������č� ��B�@_O�,��Z W}�\QQQWe�ţ�sk����ѨՈ�.�*��It���H<s��1Լs�3m`�\�ߴף�퍳u�[�t�-3T�"M-�cֻ�[N	�W�i�ik%~]=t�;�S�^��V�($����D'�E4ow�!L.�Pwõ�@�W�pn9�)s'�b#{U�IH����F��g�宂Ƞ:�24i�bF���z��O�َ����#Z{��Q�<���ȗq,C[����N����+#��"�Q�r�(��s�R�D���Od��a<���ݼ�����򽳙������1wc���8ˣ�����'��'׷&�p�닖p�(��֗2W�@�Rix�5]w�"�
l�/X��^n�[�O�ʭ^KL���������'`Re��CL�>�  95����ǀ�S��OB�$��4Ұ{�Q�<M�O�}��@��6������Om}}sGJ�k�&i�̃>_ U/�"���:���{S�S�'f���1eW��"�AuG��q�3�uA�'��}��<��,i�~�N펀mm���oOl?��`G�ҧ�I�Vj���ǽ�X�ˑ��l-Pr9ew�Vz�cs�45���5��1��L�[6�VeL�{4��v��Ę
�><�:T�D��	�Rqp��ɚ��2c�EpU�ƉJ�t�%"X��ޓf	�iWyt6�ùV6ǖW��7�ʑ�ѡ5�`�� `t����ۡǂ����m�K�x�F?��2'O���������]{��������S�>wiO��#�$�,GZ�rk�3�
.Ȣ��Ip�H��8�z�V܅x�8��P�&8���8`OޗC�6,�w)�
��k�w����M�����x;�O�a^F�j5gkcURF&��J+���c[���9�G�]�KJb݈oYtZ��/]�oұ�x�N���f`F:��C�C,r��G`sI�0E�4���>���6&$�Ez��ua�ǵwůîE�\��v�-��f.gs|�u���ͦ��)y&\ Z[D������P�}�*��������	�eIGϑ-��z��׺�	���%K�Z�>�\��2L*%��Xuw��+�BS�F�.du=#J���ȏ�����Iͤ�FM~�0g��p��?�"�]#�S:Җ��x�A�lQ����<�"�|�TW��]$p:�0+I1�S��1t�N!�C��t:�V��ká�}T��*K(�@J�(C�PC?��O�Wq�^����ժ�T��u��b����-g��7�fո]-�α�����Z��ߵ���Dj��i�o��7 � ��3NjffFa�_\= ��̛���{�t �|��#}g`��]y�����&��:Ln�1��0����J�����`R�^�1�#���ZaD,��K�dC�<cU�$:��s��t�b ����ge0R`v�>��]�!�ָ��B�g���ZuǍ;��E9k��0�����[��w|�o��o��G;�������*�/�����a�~�'�ϨEc���"f0�a�x_��Nd�z������ң׾�/��3 ��������^����&�H�m�GDv@�e9��[� �j`e�⁙�gg�P�=S 	]<������:�*ץ�|2B���@��5�����ͽ<�v���#F?�O ��1����G��S�=�m��'-u�ԭ �J�������jm�-�۽u��E?v���㧥���i�6͕����-()����Q!`��͟�(L%:�R!_���\#�WmnT�����+k'�r���,#"#�O:�ۍ�����Cuuj���jޞd&�kh(��5YvMX�|죅�� ���݇��Eͼ~�e�N�W��#�@�w��E�4Kl����ov%44t�&*m�u[B�Mu��L�@��dN4{��L�@��eFJ ��o�G����k���M�n�|}��rI����2�i�!���2Y���2e��5�T�GJ1�R�"X�߽F��u��笵�`��d�FJ��X�	*�z1T�U��EW�S؄����?t�l��f�D�v���
E�,�a�ag(p���H�x�܏��.�J�� +��j���M����;���Or�����篍��8�jS{�Z���$����T>��u�6\��k؄`{|�\�������b�}�>�`/_N��2T�j���%`��}��f����¾����!��؅��KU��8����2�:��O̥�*����ED�2!b��f֜��M�[�~�x��L����� q	����0���O]⤳��~׿;�_���wJ�\N�W���a=>e��P�eh�o�F���^/�� L��oH4P��$
�eU)!\�M%Ŕe)� �8�rt�k�?W�\Um臔���G0��ue�P�l��ٵ��Ժz��'���S�O���`񓶁��P��h�j8�����x{�-�B��i��Ձ����X׏�(S*�a���I	�E[���ź���4@�� �<Jħ<���d��|�5aD7q��Z��9����Ш{�������v3;�{��]	S�l.����?�i �r}�����|�\���m}��M�0kјwAu���s����\����V�{*��u��	N� ��6�:e).��x�sh^�Bh�s臬'�&Skp�1`o��]=y?t����y��ڻ���\��R����ܠ$�-���Y4u3^}9����U�.kL�=M`�7�ӨŃ�p}mm������Ղƾ��\\̠}����y�}��!L`�~m0�fqǕ�+H��D�-� ā~8g;�d��O���4RI�p�+q	�k��G���5nr��T�jf������:q�0SKtB��T�e�3V�>�jc<D�y���	e���{��+��B8�|�i���0V���� �u>a�v3<rU�x�R�K�h��l]�~}l#�	��+uR�+�mK������T����\��
�ٯˑ]���"�j�l�6�D����nj=i-��r1�S�G�W��fx$<���������.��33\�����
�g^Uo<P)m
�C����^I��8��N�x�����"3��
���������<�Tm�� 뜝6��A%4����
�a�2�c���+���sD�^������}�����\���q�ҷ��;���:�����U�d�N)���9������*A�O9�?g!�$z��}�/����?<6'A9�)B����:��ܼgI��9=�r��OCv$����r#;t�4(���}g,��)4I�`�"K�� L�sw"4�4y\��ql�s���?�c� ƽ�6x��D]vs�;s�n@��y���H�Htk�@/`�pW�k��UM���8��e�ԛk5��:S�z���]o�^��fO����dt�Y��=`�p�+,u���鎵�����Jh�o�p���W*auu�����5���S���`�=�ύ�Y�?����P��~5q���L#4�ҲuH��#̣�o��5��Zvf7w�EG4m/�hq�U!#��.�p&k$�è<u�ģB�6����\�ث��s�'��=w�����I��Ƙ|���ר��dY=n��d
����c�0.yM�N �r4��0��+�iM(�}�^���/�S�Ǔ�]�>3!��_�R����2��G�mʩp7s@���%�m	��Ǐ�*���^ [s뾖�	�����76��O�֌�p��G��ᆿy��{�h�~��ĭ��SUyٯ5y����P#��Ȉ�l�zD�nKCEiM#?䙊�S��.y��>��䲽I�+'��D[�\0���B��re�N�&4wT#�U��aʝwonNO���C�ﯜ%�#]������`�FR��":�XZB�4$��B^Flot?���u��x~p��}�1��oQ�b4\w�@C?	��aO�j�>��@u���]j�9g7�Rn�/�<q���KF{1K�XZ���g� �h����q��Y=ȗ�#�-�K(�<8�Y	�G����o���'�p�r��|�-T�j�����"u�'���C=k �`����(8s�$��uuE@m�s��%���ijn�Dfx;�K? z�zͰ�RH@��}u5�̹sG<�d���'��;�6~%\ztb���  S�([�Y޲��f�wn��|�Z�f.��R�� yQb��LJ��<�f��ZA! �r� m��/H�	a�e���{2�~Mg$$]Ꜣ'��Pb��P]i{�g�N��qP�K� ^�ۯ�Ox	nQ�
�������#����y�{%=��������<}`D���*�j�J�]��wf��؇��,�7/�Moe�MX��,V�ط� ���(�a(xӲ,�y0�����k+���t{�J���Li��2`��I� ��	�ښ?G�g�(U��w@;EjS���Z�<�|wJm�?#W�b��{�''m��`w)[ȳ����c��#!�jI�X�ͧ��ҁB ���y8/����N_Ҵ4�!�I	,�?�z-�M$��gp�W�V��'�}�0IBdN��ޔn����DNf5z����0C5`ڤD�2�Ż�ʧϽ��W�9}a!�tdE�s�k։a_N�@�b����9��<'!�v���Vb��Q6%˾���x�<����)�o�u��:�tE�z��k[(?	�c���I��VNĉT9��[���9f��!9�G�Z��n��^� f���9`��l����n��������V�%�W<�¹t_`> �o������'��qRe�4��p�-Dv�s�{Xuସ~��s
.��^��J��+u�VuV�_W�'���'�5r�j|FҺ>�_O��`>;S��+�4/.F��`Ѭ����e	\����\�^�:�4~���/������. ".��1D⊇K)ѩY6o}v��1�T���\��%%Ά�d���;��K��2�v�4�Փr["�i����z��W�\����l ���$�pf"`�GY�R�1恫�[���>?���9��TqeY�'#�͈z����ԉu��W C$� �s��G0���!g��V������W��:g�W��Tr��(��l{���t�H���i�Xﳿ�O�	Db�� )	��m�B����g��#~�Ԗ�1�&^��q�9���I׺���+�G3���-'����:�_�nN�-�V������1���!s��H�OdL�<� ���(W��ts��`���t��x8m����6��Ʌ��J�i�>k8;U:����^w���K�o�pj֑�޵����<���-���GSf�y�8��$��������1��d��.)h�)��y�Wjw#^�zՂ���'��K���c@U1ft��#\�\�K�i7��:;;�R�9E��>��i��n�A�4��r��bI�>@V	w� J��Y+�2b�Ļ�/��F
{��jͩ�&��6'�P�Y��n��e6H�\�x�����n�\����~��Zk�p��2����P��D<�շ�`���F�=��
�a�^�m���4��Xd�5�w�1Y��{�O�cO�W����Npq��j5�E=�S ���R^�F��6 D^��{��#b\]����]��U�/�G,|k�V����q���iAn4	󝁱����ʐ�%���K.p�w%c��J�0�����H�'$ �v��O�v�Y.�j:Y��?q8�2*Y��f�_*Y�-l�J�cV�w~���r�mk��`@k��7�ˎc�	���ؼh����.˳����1�p���
���H�AI��D�1!-
��Z��O��;�M��b�/\�Z5�t�����5d�-�KŲ�
!,����4�G%27�U�c[D�	NT�X�	ɝ��������X���5T�9�>m0yN�8Ժ�e�'�=���1©��B�w��$?e��P����Puu^U�(�H�?Q�'�O�O���(1Q�JZ>�I�;�P!���Y��,��̞�������׉��vQ�����Zm�Q}����iհ^��
�7��`�9��tx��NV�%��R'���T���
��,�R>竵LN�i~�H��lR\���t�[����vb�[o��0hr;�_*�	�|�*����*_��B�_8E���F8�$��a�){gk1;ƫ��"�}g!Mګg��;w��!%b�Ef����:�$�������8�U
n/�hXo�������8ͽ2�H@�VVW�`�*�^2B$�,Gj���l	��a����^֛��;Q�o�D� #��Tk�@g��si+Af�N�O���G��dzp�_��늄U�bT��߽!��A�'Ud�N(}�"6��%�%���R<��Q/Q��\���٘��ۭ^^X�p�wo� ��wL�~ 4K"�+ǃn�i-u}�����Ez��e��_%�%�s��
��:�=����_���w~��"eF��+�Ӯ�z^���W�����b!Wt��;b�,� +�w��ׂ��y�#Ҍf��&��� ����xt�G�()r�$��l���\��i`�D5��z@��w�gO%�vE�'&U-2�pN��vTF�Rɸ�+|0�C�Us�k��/���6)�'	'f�c�C��;^3yv~O���kA�o�
~&�r�ͮ3��[���ٻ�t��P;LtO�,�����{���p���qh�:H�+���i��9�9��v.��w�="�,���KPv�O�iZ�k(����]�z�^[����DVu,G�WV^�˿�ELo}Jgl�(o��R(f��~<`�Ԇ?�*�8�-G����w�>�/N��d0I�=ԍ�?Ƹ��g�R�9�m&� @B�%��d�s��)q�#_	VL�����TsvU�I����U��9O]Jdd��?ؖ������G���X��κ���bd��-��g6-�k �+���W:^�����Dx�4���U��k.F{R�ǂ���o˕7sN[�(�����������x�O���C��Y�Z��]_0ؙ*'<����x5����.��}D���Ȋ,7
"8 h73]��S�4�'e���|������B��~�\e"t���N��UŮEF��$&Z@z�·YN���cU�'���k��0�;�b�u�Ⱥ;\# �Uc�hj���/������4�ۗ
�f�N�<�U�,o�6yThU�bu���Ⱥ��Y�q,1��^�Y���4*�eo����I��?��i��8�������A���>l�H�[�˔DGm�;m�	)�>�Ymf��}3��F��~Q�߅L	�����
H3q���M����v��Y�~�ԃ���h�f�3��#��U>��H��z��w�եjXWq�8�Г���`�R�{��F`���6!�����_<���t_��]tI��A�d-&C�:ˑLHi��y{(���5$g���M>�0E>��f�����,K����f{|c$3��
̆��C��ٯ�T0vӿ�N
��D�zpKj�N�!ჱ
�xdm~{!�@�-4�c��o D�����y����j�*�`�		3�-d���J��
��>m,gϣy����jc2��q�
�ATB���F�k�/�J������#At��6��Iʻ8v6��<%1����sR��ATzЖOgC�Qe%�g��}�ޞl<ԟ���$V*���m�9E��|�Afшx���sv����4�F����y�8�K���B�n!�-! ����롅ٞX��85�*~�����[J�(�ߡ��������_U>�~�ֶ��S�����즋B�aM�j����eH�E~�G���s�Ӂ�.hᏊV�g(�R�4�̚�L����a���'�ș�0,ib��8��j��L�p�� ��P��Y� ��5�M�svNIz����s4���1&���6�Wrk��Q��u:ܥſ0yV�_��[�v�f�����U����29���eCť��a0Z��7Fn��l�ѵ�k�1{��� l�~/�+%@�Z�>0R��+���G���ꀁR�|>����Y��Pmio�e�	f�
�͛+�揾W0��ͤJ	�Cs<mG�|�.�XTʾڑ�"t��~Yg����=:�+�v�Z�}f>VJ䗢?���/�|�t:���H=����&�8RS�V\�U�<~�|H�d�S�����_l�b��Y���9��'�����0u�Pu�'��D�R!���d��"�W�i�,���nJ�%�(�i,[��6d�ƒ4��6�GR�s=�������l��9�����:�Ϲ� [�N�GЬr�h-�;�����
#gB�)t�{��BY�Y���e$��،�	c'~-Z��)��S�����w.��x@!�o1"{K��G�m8�B��g��R���b�)|����GU�dI��-��>_���[ɸ.�b;�G�Mْ���2Ic=r�dť���zd6�j��*?��H ��m�D^�2�_<�)�<���d������x��2I@)��~��?]n7���Kc-�ݦ95L�� }��]�WF�����&BO�*�8���VVƸ��Eu�GV�b�����:'{(	ۍ^86R����W���{��Qv���k46-uf=ܨ�y��8ӡ9H:���eڿڵy�z��$�!����y��@��D6t	���ESjW�;���&'שּׁ���U���}�������ǭ��g}��!׷qQa��y��Q�����������Q{rҬ3H�����9]epÍ/�ԍ΁&+FG���ߍ��+R���k�5&j�b ݅3|~ɒ&;v�9Bn	c�#|�Q���3�⾎�u�e&�����'2(��)4u�wU���_��� A������w���c��̅�Lc�G�λ߳�8s���\�쯌������rV�B�PJ��ϟW���o�6��X^�ʾ�:���q.�~%(�J�GFF1�a�7�e�-�A��	��7.�v'��̦�c��� �y�w_�d*�K��-��P&�0�O�Bb�'1�|�M�"#��{���!Z�c��l��}r�ʐ�k^m���+��
GE~�s+'^�:R�9�����OY�F������zq���:�*�Z��W};�x����xܕ��צ�k�iO��fU����.1�	Ү��+�z�iL�ܚ9�B��9g�4f~ ��e�w��'w������������B�������9DIT���J�E���)������Q��;�)�Nk�Ĥ�Z>�y y=CI��p�ޯ�py�I�lRS�C�T;�W��^K�ձ�j����ih�ÝJB����CU�f�N�,�]
l�n�DR�2i|�7*����)�i*@4���AoOb�s���u�G4:F�ħ�n�U���Q������r��4w{���c�";�qʠ��{&���z�Ev��"_S����5%"�V�����RY�s�$S���)���2�=K����Guv�JJ,����7E�����t֊�sj������3�S�k��9��F��y/NI�K�������� (�Zg�s95H�XG�˰煈�b2�a�<bp}�5��u������%�9�mz�4P�%���4� ����KN�M��br��xZ;������;,�T���qB��%1��Hw���	oE�:��'�i��ΰ��O&OO^L����F���V�ĩ���.��yk'˖#.\�����lJI�\���h  rYv��N6��fw'u��������@�^����R�a1_���1�'���=�������4F_^��n��������&��r��WJn���i�Ѯ����e�;㌻YB���ˬ�XSx�T��O�=��J�ӳ��u��Kn	�3���\�̓� *��R���u��q'dE�:Ԯdȃ���}u�qȣYKZ�ȃ#~գur��"�2�.�c'�.�z�x���y��*�!F!���ڽo��^,�`��j�9q�&o=�lI���e������kR��%���)�* H�qW�pxD���'Y;R�'R0��!�.� Hj��1[!�5Ќ�G��샻��rf�d�_���2����3N.#��y'<������W\�XA�:��K�-��bY�%�cX�HF<G��֟F�jX���_U��T|�}}�;��6摏ww���&v[˱�$�6�C"O!<K^�[,��:ܛj��5�pZ	���7�|�]H-S/��Y�r]c���S8��Q�hz;�%�P͠_���;��:X/�dԩO\��_Ə`}RKV|��
�H3Z�Sg���DJ�`wIO͋�s��, �+X�w:j^���2�Ǣhl���!�c�I�
L�֐V��>��Sןx�X �t�4m�ⱡs1>6�LC��y���D�?П�)�����JcR���-Q'Ǒ�7�����EE�����fy����7G����W\B�E�Y�,��@��N~o
g}Ib��Y���xeͭ}�|lN���ӑdR�1�j���3w��-m8�:���y��;ʟڭ��黯�K1wL�r�CsPq_�jU6�j\���p 6�9:�9�ů���܇��� H���s@#�cd2�L�x�8r4�xc���]�qu��s;J��SkK�J}�P�!W=�S
� ��W}��I:����c��<�7�5�o�e�d�&�i˷=�����ƛKg�\���o� c�ϯ\���fy����5�Z[�8�+�E���1�]�W}�0�/��	x����h�72O|d�S˛���>�3���ۺĆ�c��Z�<jt��7����a](��Xݜ!ɀ�hA��i��1cy�.�#&&��B3%Z�4	G���r�z��EC ����49%ǒ�~�M�'=�����*V�����F�� s�p>|#�Q��^p��Yg�~������}K{����Sa�Bj�Yݗ�b���RO���{7Q=}���)Aɳ:�Q6[�|���'5��o��i��� ����7Аw���wR�_�����}TK,&q^S�!Ü��9pES�%M�< 'PS�����>��/�v��0�YǷ�},���QG^��cRD��n�T�(�g�( =#AX�Q��|��U��Z�|�
��]}'݄ލ��x���M�:��io5P�𹲗�g��d��� w0��M� G��U3��ǥ���){��ñd�s(�zʹ'^ ��BO��0�X,D���i5���绶��GA�P��m+�u�m���N�`u�9��]�t!�]�L)G�_0]Q!_}��1tW�)H8l�jʣ�d���L��P���H܉��'���=/ZC�~�i���1�?<�,&�V�[��'��Q������=�j��,�:�"U�/��޳�5J1��� 	~U��;�2����Ȇt�H����;s��D�_޵J��B��@R{�Q�d�y�) 3���I,���< p����nk�Gjʔ(��M�O�$�*�cȐ!��H�`�%�T-��D��y(S��sS�K�hV	��%��ЋA�־�-���U{�?��*n�簩I!���[�ISj�/2�umrk��L��<6��︨ޭM��w�ٗ��ř��V��B[��a���dJX���/c�\��ȩ}1�=���d��[S裓y�©��'yIƕ<{����I������`My:��*tAK�2�$�U�(�[��@�O�i
�uN|�-a&.^w�;uZ�Ur����T�0�6�pI�vU2:\:%�����dڶ���v�t2R�q@��y���{@���lиXL/kG>:+�Ur�>(t�-+����1Ш��KT'u]�nO�!_b�;�*d�B  /7'��LJ���ʚ^�=�ah�r2��8�7�졲�;� BD8��HT�I���u ��e@��H��+�u�2��9��`��Z��Ȗ�e�҆�wS�a'�dƢ޿� �Z^�θ�iӵ��v����mQ�Y{��%Q2.j�|#��	��.�Qz�W����41�:#H�9�S�E|������ڰS�U+��1��)(T�%K
�Y��Hc1�-Uf�@=Fq��&R,��_vwk�"���H���j�����GF�_�#���v�������dN���y�h��v8��_U3ڿ�/rn��z6���
�8�!U_Ѧ*G�7��df	�\^�4�%*?�X�[�Mv<Q��xE����r'o\�ԥa����q�b�K54��U�.ego9�L�Nc�b�m/�V9_����hHh�=�����~���0?$�bI�3y���aZ�o�%�,n�#i�oڊ��3���9��RI�[m��:hAKO�=�EĎ2���~EN��v�X������x�r��C�F��Ɔ_?��*t~o/Z������wW�x�PeC�a+����m�X�T��OR9�!@�U�W ��&jF �N&~Vm����tH1�"B:��Z�	�Hg-�8�P5�Xkٻ��Y~�;�ˍ�O�(�U,��:{ǋ����!>��g(FE����c�U��wWtZ�wt��ך��O�=����*/ k��͋d��pAJK9{U1 �͔�z�GGd�:�8�'�8׵X3�3]D4��Y�_0��N�����^�����x�ġ#P�]�Y�s�7��	�,���k�#�}�I8���w�'^`[9Zog�^���Y
z��	���rm2�u-'DҀ��OY�J�F\�;E�<u`���h|���`V����b��Vd�$E��5���MB��8.����~/�i�C���v�����L��j���2�$��g)Y,.���Q���Еgr,����k*�?�,���-�4K'itP��F�3���������V@U�lrv�꾠W�� <ƍ{��B����Z���k�b�\ƹ����eu*d#I8���L�Ŧ�c(�����!޴��*�3��ȷմ�_�$��6gY��$�Ϋ�ǝ%��?��I�boB!u��
����ne�`��C_H��R|�m�vm?��!}ڵ�[�c'MqϞG{^Dd�w	�Q(�FҔ���)�=y�m�5��(a<� .�������	HD0ż͐E�W�`s�Fɱ��R}��f��qT�hq.����A�Z��u�wG�<�0��iTv�̫��3��R����Ω� �ǯ:+	3����"|��=�`���`��j'8$�� �Ԓ�A������GR�*oX'ʢc�����e�����>��!� �������aC��|�2 '�(lx}sÿ2�V^����Eؓ����q_���4�V�����T[�|�*6uZAɦ��C�t�.@�Y�L:;�zx�����w� ���V@�v���ax�S�eS�P�K򤰜YjQ>���ePGx�]\򾯲)�W���Iꝺ�a1��<��
8�p ���ä�>ÿV�J2�!��j2�!�)P5FB%��J�:��<�2vo��ku��Y��Pio��i���C�O����>�v�lJ�c^m�� c Һe)�-�"Ů�@ڳ��CG�u4���G߂}���/��ۯi��b��m3]Z	:h풧+��#~��ΦUpc �J�(����M-���L����
�o�[0�2�`���:��(-���+%��#s��eB7.���w�.Ze�޸����ikO�.z�I�toj��/,�>M�r�-U����GrN2{� �������^���*$����f����o/�V>>d
L�i(0;@lH*����,�"J5���cQH4ܝ>d����3*��V+�a���{��4�S3��g���^�?�ݯV3N�fu�Sdc�_5��'�ʰ+8(o�>���3U�5R{����Թ����sk�wl��S����>�X��{�X����!�-�0�� n�6�q�Pٻ��L�"Cf����z��7�����HGs_������`B�d��]f��]��b?�Om>�T��l��ԉ*��[�&�YW� .{蛙������}�e��y����q��V7�f5Zm���Jܛ��|�Ϻ��O3o	��U\��3f�/3��/���
f�/�/����C���/��'vۘ�K�d��Zf<nME�DweZ9̗7S���)B����)��)E�[7�9	��E�P�˄���:�$RI�M,�s���<K�0�����r�F\s�I���C;�_8w	l@� k�J4ָ�>�M^���B��m&�	K����|�ϸa,r�շ'�;���s+]/�%L��d�(c:!� ��?II�nƸ��$�/斒Z����d�� @�ewX3o��ť�a�`]:;M�<�5�<��� �ҽ�i�݋:E3OC���H�"aZ癘K8�����v�ޔjp����E�wc��]�ȵS-c|���dV�Q("���p�s)#	��'��\����%DW�K��|%�ibκ{�U�﫾K�Ctk#�ӄ�4fw<��4QZ�;#����:�zbq%/:�*"	qB\;����-��1e�锓��]+�8e��]m�GMժt����� ZvO�.�qVhM�9��ЅoP=]�L��� ���k���4(��?�n!@�W��!ŗ"�l-�M�}��Er��H{WOM��S�A��F��*b>�t�j�Hq"���I��xP���sSu!�P�qI�18��8u�XPl��$�yM�K�u���w�d'C�J3�2U�Z��X��;����[���ӗ���#��mS�4��`.�WFP) �3���:�3]a��1�C=��X.�!̃��v��7�֯���F�� �6c�d���|�8S��2�x��r��'� ��1ٝ�K%�RU���.�u�i�W��Nۺm�2�f��q�_�sk�y�S~ʀ�����D�l�|A��ޜU���J�R��=K�@���;fW] �1d�(��CZqz�!Gx=�0 nw���1@.�:��a`8|nC�7���n�)�8U�9�Ԑ_���m��#�B��W7mAod3���g��� �d�ӭ��[�~��-�(x>ܨ�p.�3Ic�de��8=p��ҙ �R�t2O��J���>�'ט�zJ���sU��`�4�Ql[C���`J���w�����C_t��e�l�E��+Ů.!'>~DLզ͠�4�z5�� ���x�j&h��
N�h#�m}W���H���6{ g
��G�������3- �ؘ�6�/������I# �D^��z-q7J�vC��(��|ۼ|6����'=�}'Ȟٵ�����@�#��;��J��N�Ψ�Q=/z<�����O��/�!} �J�P셠s�v|�W�Kڅm͟~Ff��Ev
��C�n��#��ۭ�/�Z���¤�'Zc�o�����`����
����^:Zq����^br_z%u�WQ:�l�s)�f'eJ�9VI�ӵ���S����q�K������?�*Q����Im�����k��p��w7j*B�ұ�(���!~�G��v*���r�"�����������5�m���j��3��-ô�@��p����a�y�+ɜA�K�������	]:��̮&�rÜ�*�� ���G��&��� �9��e��6�R��L臏o�8.Q�R�M��"L|�]�J���y��G�5}%��>Ⓞ�g��z!��Y�e[ ���yM��ݯ31�g�<��mL/#(�W������Lq�j���3�5z�i� ���^KzǍ��!�MC�I|C�R�Đc�1��9����ڌY���tPS�'��B�C���k .���76�+:�]	z遤����� �LO�$*�-�|��n�i����
�7:+��{��K;�2����SX��Z=+84���nne��,�bl���ş�C�\]u&�tZ����>�݆�?�-ϋ�g�e��ͫ<���d<��:����/|����
��v��*0";��Pť֮�!D5hM�����* x�Jg�:��9�����F�=�}�Y$�B]�(�k
�o��PI�9y��V����[Ex�/:���3[�cT��|J������$G�;1�����/��@�ƀ>��Jd��K1}�U�.�W ��&��s�Γ`H�x�i9�f;�\�Y8ӕf�<u���l��	*'�)Z%�B�8�ߣ�ݏ.�Tx���5�ǘڜ��,+CY��c,�/Jp�N���r�-��7��VOb�5e�S�[O�Ɨ��~-)����i��)s�P"���&n���s3S �iC�R��զ~����_2�ƐZ��|����d�&n�?�^��X�\��{���Ǚ�k6"�>@ɔ{D��?�I�āp�W�&h��XL}�sJ·��M��"�����An����U��=��Z��!��WU<"�V�ږ��c����x�G��gE��|#
�|!��{����~���뵤�O�yCX�`��̦�}/�Z'���"�$u-�I	�jn@���VL�d���[��q��/0L��h�{�ȁzV��g�n�Kťa¶���t�$��[;=�\�qח��gY=:w��� �J���E�_�V����}��Xl��>���SX}�Q�u�wA���0[��𔏾.��V�ǫ�<-0ܮ�]����=���9!l)��S�N���J�o�[W��朐�aNՍ�vZ�#&�F�xA���,ɱ���]=*뒪ő�J>��: ����Tu|��9q���`��lċ��>�,�~1
)�K�������֎y�)�S�N}�"N1R�rfi#ūzٟp��@���[��[��®��+k�L��;
�0�[a�m��=���1R��� �v:_��2���Hf�Ի������l�[*j�r7#�c� Zֶg���Sf��[�`<���Î����ij+w�/=��l.�"�u�2�_L��M���L�	~�����sx�~ϵ[��ۆ�Q��Q��
�����7y�x/d�nxR}�>��5��ߖ���WѴ׃ԀnIB�������k(g�w���ʝ.��Xۘ��8�en���y���*��#K����wɳ`G^�T�U3��K�I�S��/���6rhor��?1�EJ����KY||���ÜS���G:���f��隝t�$�u(/�֖²��G��r��}Վkn�N����
�Nl����� o�Y[�M����O/�}[k8�6��kq��N'x^>v/�G������ȷ���8&�U��
'KW".�CUi
 ����'˟�,KO�=9h�x������>�w^���ބ|�
�>�w�z63��СHr1Dނ�O���g����5ӾAJ�-�a�`�-Цa��z���������?k�eKQ�&��?�7#��||�Q2����zʗ��l���4�@R|�`}ҕZ��G�񸬄��I��G�.�[��z�O+MI��R͛/a�MA�(f�P�����Z�����3��/�0��جv)r[J�����������B��P�L!v�߬���"|7��`��k����>uU��1E�t�ײ8!�K����~�t�
]��ʩn�X`�)���(t����% ��1���B��?�m|�o�K�i����Y����3	6�\_���5���*�;�v�i)���JzZ�vN��c���t�[C��h�aj;�r�����|�O�� �`��t[6�Jy�<�ZE���$�\=�I���;"r��{�fW���ܣ$Z��O4�j,?���Pz��Qޝ-;�ga���q[�fȾ��.͜k���BX<��}w>��&�2���5?K��7�h����t��]�>D��r? T.�Q��SJy�AY8b����#��S�TDTĹ��_+�@��ѻK��z�Sk���OB�ܭ]� �"c& ���Pv� �Ũ{�	����	ӕ\�
�����r�<�o�{�4�mI�93�,�b�,�� �߸?���Q�5J0d��ÂW�� 8NP���i�؇�۾��,T�F<N-g�����:nB>���-x6v��E/��-`T�d�	��8����*��:���\`�}ʕA��ȡ�r���~=���	K'���XՖ���8�E!Xtw(��5�q�4�����|L� ������Xz��Ɏ�^�-�8=M��N@��^����P`vN����W�� !�	�����l7�,cd"� �$��Wa���=��e�n)�����A��<Qn�vӘ~ӍAu��,i2^¬MF�t�%��B�@���3:���-���f�s���,�F�N�q|��v��M4�|er
hJb9����2ej��lDک�������9k�ጦ0�+�Tg�(�x�͹�<%���WC~J��4m�h<�}�8+�<פy������܉�	&QQd��*!�U�� B_�M�-K��ݹ |~�6��>�����s�5GO�ޫ������#���~ML�<�K�����H����`�+�,�\�絯�����;d5
������{�D,���T����Zr%���z���zG���ϟ��W}�n�0�wr�w���'{6��&g@�fP���_Gd���ܴ^�}��������)�`��l'��Ѹ^������a����!"
�j�Ց�W�vV:Vj��
'�8!.���0�D�T�f�3y?�L��kF�uu�fh�3��W��0`#�pB*<ʶ7Ry�A\^��#eo#8�n����#?_W����v�q�V1'گV����?�|% ue,W�"G
2ٱ������(���]��u�_
I$^���R��W��q�����*��J�mC M>Ɛ8�a���hy�} ����B���_�������Wf��ͮ5|"^M�/��;&W��вh]Z#�
b�Z�^�`�I��eNX	��߾Q���sS��/��v����f��j���a6Rf �HyA� �\1��D�(���"����:f<�`����"i"��^e�	]A��^�0Lq�X����2�RO��t�bk�+
�ys��۪���!��0�����!�%������ʊN�y?�
P�D�����}�IA62��LtV"n^��S�Z�(����(M:k%S�:�z�&}ok~D~0�j���w��.�°V��h/��x=�;q6c�"&<�*����߬k
ɦĞ����_�����i1��`�_'�`�r�tM!��[��3Xe�\��#��PzAD��g�i�ݻ�̌:�,��ЍTm�oTh�-u0Ro{jm�,3hxA�	��4�������#�������\UM�{o��!�K�d�8JR<N��%����ԡfJd��G��#�0��x�L�8����!���d�������Vn���#U���w���p�k,\����hb�=�z���~���S{��U!���O�Bx9V��c�uN�yh��'�)������О:�5D��.w��h;N��8�j�cUsP�7��D������
��߆���a��u�F��ᭇx�l@��e)�O*V;o�Ǚ�.U�K�����j��Ǻ�4�\o�f�)�����>��I&#���)ǒV�r���ә7%�U�����S���j¥P�9�Z���������]Nf��:��[m����FDv�#b�qU�ȉ����g4#$���Q��:���=�i3^�Q�`vow�t�;��E|0�W�13u�< jq*z�ۡ�<�ұ��zHcj}���X0��^�(> ��Ҍԭ�� �I:A����]�c�Yg_��>���x�+�X�	|i�<�M��U9U
/�<]6`��W����R���F�����ڿ}s��	g��,x���IflT(�ǳ*�uP����Y%\;}H���i,��m���v����{[��Q򬥷J��Y$=`������O��K;4�/"��fW���M�>�cj5|��k@7SW9C �3���_�i��l6����<T�F9�q�+q/[3'�hf�gFB��!�U[��RSy���䨡�.YvN���f|_u��8<��a���e��m�<�B�ɟHi���F	���i3�՗�lq|�f�|PN�������7��2����?h^�܃r� �>�{ԶՉ��g�zئ�~��eiO���ɯ��@�YثA��[���HYʤ�}S���o�9�¡;�N˸��s�Sz�|�:C�i���a�x9U}c�ט��p	��]������]��G@ ���-��KKɤ+�nm����E�0���E�:?|	;p��*sԘ$�q�;D;���Mԍ<���͹�*V�D��yvP9�����o0sV]����S����mO��j��\��{���X�p��u�~���5eee'�%s&�8��ಔo;�S��^Ijy�߆!����� �L����ƐZ�� J�G���ќџ/Gφ]0Nn7�N��f\(>���wo��4�����tQ�R���N�\�{�Wӡ(�y�)�Մa��P:��S��'��;��,t�3�U�3�FQ�?`^g�o6���on��1�Ϗ�胇{m���5�74��o��� oV����p˼��T-��>�������&(�Յ���v>_)���=pvE��n7��k�H��]�l�k0i\g4Zo ����b��N��e\��8��N/�g>T�|�y�KI��9�e�Z���_�N<�OSfN�G��ۘ��_�9��KPQ癷�Teԩ����T�V� �S�2�3��;�O��9�>�&1>���{z�֗�M������p���+K4PL1�聭������wQ%y���P��<a�wA]bP'��Ϊ	�ȉ������ڈ�z��������E^��(I4ފ��Π�CA�۠ 	�O�� s5N0�,th�{�)�$��&���*b�#)��G�Œ�ti�'s��x
��JF]��Q,cu/����%	S�cQ��w����a�d6ɢ���� �ր�B3�g�籆�$-��aYڎǪt	��}�mS�N�Ip�a�)ߏ*�ƤN�a?��v�������08U����A��w*�9�j��ob�{���q�	2y�Y���̓�z4@!)���3�s��^c23�Z�f�y-N(��K�R��:����2�%z������$ ��gV��/�,�P� ]ڌ�Z&q�����+���lw��l���t�6������N��a�L���ޞ���S�g��[ݷT#�'6unǍo�C8�<�~�I����$��e
^ƪ���H��SO�Q�HA���������"�����s���!�:m�� }���c&Q��� a�s�@�Q��[���pE,!ɼN@�x�Z8�z��,�U����?m��B|�4���6Qt,�wn���e�1��W��}m&!��������S��^������H;% �.=��40/�ok�vp�m��)���Ee��^p+� �V9�iSBp�@4w
g>�J�*��ix�8?q_��z$������E��;5���W͘o�e:FFn�!$���F��y�^��[� ���yn�j���_��p6�C����L�;pA߁�����_wಾ+��/��ή�S���b���G�G�\�!�_����6( xߡ��FA~Q�I��?��t���X�#2�p���sܫqT��0���#Թ5��/�V���xr������O��z�JG�JB�k��8�Y��Un,(S�����q�>�Q�׷�W_v��҅�Wmv]����p�����~7��n���k���UNH�[kD��=�W[���#�̢�p�@�u��qׅp}��F����^��w��E�hJ9��<�W9Βp��amy=j(r⥥^6�Ҕ�R�^Џ^���6x�Y%k9�vfyx����>���R�(������8b���
 $�;�ı��q�V���
N3�Ő�D��������0�@�*��Z���-�V��!"�)�u�3�̬��<Lb�(����= �����4r�E�������B��[���2-@�6�c�>;��p_�;�����o�:���$[H�k�-<K���
��<��)S�3�^ʀr�8��љaL�f�G �p��-L͜CT���'q�a�k��q������ ���Q@��m$8��$����5�ʔe�F��Y�`�~��q�㭉a���8�K�X�&�2-ӗ����3:�������I���o�Q�P��g��^i�,�1��͍��-����5��51!�A~WM�c�t�pteS�F�&$�5z�=���F=�^�m�U��\ރ�Y6�&���p��b�U�H�����H������er&�����00�w��b2��PX� ���e��yDb�E}ݨ����.�b�7pdW
�fd�\�\�~�7���3�TJ��$j��7:+��$�庞Cu�Q��Ҫ;  ��̐���	m���4��7��Ϟ�1�̈q�{K}+~��wT���=ۈ��U�n!�b���,_1��{Jl��U�~X�Q/'om���M�LmE����~�mL�n��O�洄g]����U�s�X3��	�df�w]���Elt���]�V
J��Hܢ�W��jq��G6���Z�Cj�U��g)�3@"Rݒ�� yڬ����|c;/k톸'�uh���1�p�N'��7jL���������O����tQ_>2@N�NN���*]=�Q���&l7���+O�� �\Ad9�z��� �����@y�@�	-+�g6��I����PR�&���LI!���!�9��)����gއ�E~��H[6R,����籲)��p 庥˚K���fVZ����/�6��&��
��܃C���dn�> ���o�h�s�C���h��5bdddڰm�u��ĳi�,u~���9�M §S��S
�����Rb�j�g�^��L��R�_T�^��/�j��d�$^_��4L+��܂j�'3a$��;�T���эF��i߁�����6w2R˾��c��S�4���u������#��k{:�4�p�5>HKc����s��EG�M�4q8"�qƞêW��o��z"&�]#�o�
c��h����Ġ��P�Wy��_Aj�4���$�p�={�a#�w����w�#���R���W�lK\��U�����d�yM�r"~ZG�t� ��\��m�����_�7�^b=�;,K4��oߩ(����=�NE.J��"}�V�& �����<�[+8�g��?�=[�T��y�� t�ν`p([j򽜐�$��B[-Θ^�>[6��	�v�[[�E��a�T�RJ�<��ob�[�r�M�5�.ne�~���u]���b�i,�V?r��E��n�pM鱙Rc�]'�V�p�k8�����|)�z�ӮT3��zX�z��I�6Ψۀ��L�7O�n����oܸ��?"	I]������-����nϯ������Ks?_˿�ib����i������ϯI�z��#�Oal�j*}K��w)	m���7S��ۚ�>�7;�R��4=�j���*�BŤr�޷<R~���T�Yf��Ɏq����CG����t�R\�Y�	�蘂�~��.���%��(�X�����}�Y���Yb�AЋ�Ft�������C؞���9��bJ��F��f�{6欮��}�7Ͻ����/J��je�c�Fv���S��z����^^%dH��#��n�j����F>�Jh�wH:#z�	 ���"�পc!3B�5�#�0���vp�_#�?�y<d����$S��xR'�������{�7v����s�U#�OB���s�kz��D�r� Zg�C&8��_(�|��Bk��
��j95+DMo,_�� ����h
����JY���]Zp��/\
?2I��h�U@��o�����n(G�����ұ�8��k���TDW�ܝ*aw��Y�Idn%&��җ5%2L�������_S�_�~:.h�^�uM�ה�pXiBR�>;��G�O��2{���k��KFE���5���vDP(���^�]�s�*8}k��F}����	����}#�*��`w�8w�(��7�U�b�3�T?�n@���w^�����{ l��z����!���F�,p�{��qC��0҄>�?H��@����;�X�Q� ������j;�O�:�H��SQ�J��utAmr׉��V�n�P�g�Q3#t>(����a1X�P�p� �`���:N1C���SU�Q,���)EW�8����V���%D9.z�Mk�1�+ں!�!۽�6��$��),����d���9b[���	Z3U><O�R֒�Ch����s��,�7/��������aj
�<h�׆�g������F9w�ޭpy9Ŭu���k�4����-�k�eS�ت=ے����]a�gHmc:j�\�ӎ��$Dr;0;�%��8�ǛYE�-buz2�_mYwkQZ���>�����@v����e����sV�a7
`��Y8�l	��LF��(
�vGoe�T6JR �ŗ�t�<Yq�ƔR�4`3*����-����� �)�S��*^����x�g�T�t�ʭ��l�p��*�m�X�4R�O(pF�;����49n3�ޤZ��qQ�v���}��?�O��E�����#X}y	��CZ���>�4wxY�2��n�r\�Ù}�J�5��ea�w��8��"N>�m�S���/�E�3����Uj'�C��,_�Ip�;-w�����A�}4"T�v��!�-`��y'����oc��-��oV����ʄ9ǫp�z����Ҧ@�d�k�[�K�������J6����[r�,#�&�W~��0����ޏ�J2c�!V����ŭq�`�MI��y�.s,>K$m���%9��k�׉j�a�3N�5��	�[?��@)@������P�ޟ������Ld�p�If����dh�����y���:�x�ؽ�������tZ�m�E$����#5��5����X/ n���}�����e��*��l�nm$��L�B�qR*zK5�/9�DaZ��{��$��W�۞'�˳�r�d�!����~(H�=�&H�X�����&	��^2��V��p����wq�^b'�3��2
��Ug^;�8y6��}]M2N:����5��p|@Mu�Ϻ)�fH9���54��Aڅm>���|���y6�R����pC�0�KunZ�_I��.�p����������|����Eb�#\f��3��ц��I�j�+B�Ƥ@�S���&���!�<��/XĶ�Yg�G{i5N$ܨ�CC��gb����y����T~d�b$�h���?�1?�ɨ�ۇv�!7�}���xAS?̼�*��%�E��n��11��L��o��(���(G���`���e������ m����&�]�Q/�A{))�ŝ�����$VNN���R"�Σ��Bud�%Z�)w���m���N�펿���/���_(C��]���uhf9�B�NS/C{�d�����#�a�6': :q�9xu��%�5G��%l�έ͇�� _A�����(J����4�Q�iA�Y�{���2|���SZD��zb�� u�r=���#Qt�A�@��c_8܅�=�Z�7������c���r��YT�x
�k<�c�sIS!�"��~8�(;S(>_VgKt����|}&hT�MwI���l�$14�-hr�5ϾƘ��xH��ϒiwU����/�&jǝN���.Z8�������1#�*o-\���P�{Tv{����	��8R�Ў�*̶d��	x�S0�'M�>�U� �z�������䮋��K��=Nm͘�K%��L�А�����W�+ޭDa�O���P3~@�Y���7���������)K�-�GaDvBB�lY&e�w�,�}I�(kJ�oI�a&d�ƒe�K����z�>�?~�[��f�3s��y]�<���<������.�zE����uL��J� Np���u���k���s ��J%�ˇ�}}�f�Y䦆&��vI�5�2�Y�Ҷp�d��ᒁBMU�4���>V6r�Z
v�x��6����{���Nt@א������6��T���֩�Ï凗2��qK>^���:e�����Uq�M��t�`�:B�Z�9�a���y�|h���u��q�M^p��8��,T����_�޹T��ݭ@x,�Ā��\��Z\�>�j{���g/E�qO����p��:��ZQ(��$!�x��lmm�(勵L^����yc0���x�K#!v+*��¯ߢ�)u���1k��� w+�@�����N�	�J���u@��E��!�a�SV�Ph��K��Zp����eqp�L���n�\���xP(��>&v���n���:z����������n�_]~�?wY{'_�vZé1�z�
_*��`��k��P�|���P0$|�]��q6�܂¼�k,P�ؒJ�t�� ���[�vv�b�_���,�l�����=��)Of������ݟ�#�g�45�DJ��x���ހn��q�m�?��J��_��z�ޏ+.��8�36��o�ɫ�,�7p��ྎ0��+���!]O��W�b�h$JuzW�L��� ��A��
����S�����7?Ό�|w�.!y�����V%��h�ھ_�	����g���衰y�L(cԌ�<�_[iii��"�R�����U��f,��� ��S�f�EnB�R�ǣ�5��q�0)2Lq�/�n�Ko����k�maK�h+p�,Z6m���hc���=���p�b�O���kT1�c��ePӘfM0���蝆,ߎ�]�P����r�-aE�r�W���a�^��3��u��#����n6wf��
����)�Y��#G z�F�߷:��*���jX��b1i�L�pX������3���C���W��L3IFe�HTi�
�PU���a%���xr��p���yr7�d�=ؕ_PX���� �\
��ү��W��癊LTՍ���wC�P�QH��薹GћhT��7=5����jz`��!x}�؄Yk/�*a�s1Ҹ����
�0��Ƞ�/�-k��~h�D����i ���hKp�J�Rc�IH��$��%���?�?�ap3i�X�H��y4g���:0�v�/  �ۖ�� ��}+Q�e�N2��+��W_h	emb�.-�R+�5�l����k;h#m�2���$��2pa�,��=����/�M��ĺ�v�E7Ub8��A����"��v|FLǂ��`g������c�.di�%`������새?��2���F�������%��p@�4p��PA8��o���j�7|�.�2b���d��lL�v|������#b4���D ��2fb*-Q�*P�V��_�섿ͤ[������mꉵj��5(�t�6U;Q y�sYA��7�pS���@�
�2� ~ �h+	4*��1�؃bI3;�۲�]�n�����R���e勚<��L�)~dz_[؄�}��\��tC��������8�͑n�����ݍ^^��,���� r�J�Vm$�G"���8���/r��i�O�<�<��?@n�w&;�e���C����C��Hw�+�}�����؋(��`�O���4L��WJGU��N��F)��w���/蝆6��C��ӛk=��{�����ɏ��?����9u7����T���ZEJ�w C����ևE�b �V�"�U:o��W��݀����,���e���
=]���G`/Ώ����fY��zq�XM�-��ǿc�d�X��y�]�.�Aſ�2�Fq<��5� Dm������6�=�4Js�O�W�"��C�6�G˴�bi'�}��/�f�d:�eu���e���A/�/VRw<�6ݖ$���Js��q���Ѥ�8��3��,ۈR@���������7W�GD'�=���V��9�#D'�c�n����8��O�[���>G��u2����chx�k�5�87#��U�w�4=x+|�up�V{�0n<�L��Yn���h���0�3���5r2�f��V�=�P	�%���\K�����Kl]�bO^λ����0�����O!�/@{�U7�1����Z�Rp��hcС��y,��wkʂ�"$δ�N����޾o�w�nI�n���/��HA�G~0g��?8�y�t,� �2����T�C�2A�F[;����^�w�w�<C��p�p�<u(�Gz�Z��v�Vn�D�W#��x��6LvTN�@�j�)��H(%.�3ݕš������2�Y9:�v���p(�l?D	i�=Ml�v�#_|�:<�6
�텙x�;Ner�����޻�$-Ճߎw�g���m٩Î�2/tat8K�~-B}1�2Uq�S^^��/c���C}��!��Z���Y3��vqkr�V)r.�f�Ur&����vW�l��a�WSsU��E��
 ���`���e:����Uw�Y
�7�W�Xݟ@�����;�Jf�Ź��9 `�=p��(WVs��7yo�1u���8ZKp)�<���/�'���&TO$EP
X��3+�
�A����ڌ����S��Hh[�T1���9��'�n 	�( @L�j�����Q/T�_Gm��eM��o��(����ɟ/��בR�]��;������ŅE�ޢ��_�c�������)]v�6�~�P�92̌Bc�C=�O*�4�Ԅ�Q���+���{(�N�@ף.x)#�[�|]|g�x�J�Ӽ�ᡬ	+������nq�=�YGg�u�3���_�OP�����P��ip�׽���fj���u��n�eH��!\n�/�c��>*|�Χ���ow�XG+�{�z59ϯ�����#�,N��t�u��:HmF춞£z���X������E͎�߇��n�����mn��=��n½��"���ψKᰋk�`d*�N0���܁�^^��f.�kf�JII�{�F�W??)���X��p��&�{eF����C�a}�1�&b-)�6�"?�3���C�~C�sO�xE���V뻩�U�� ���Ha����I>ژ�%����mvtD�?<2���Zh���;N*]?$³���Po�<��K5������he����������o�����^w��T�>|��H�)ix��{��BB�#���k�{�=*`쨥Df�c`���	+C�zgP���7���R�Z�q,v��r$�&�����/����/�k�b�o�Y5_�m^2���xi���^��4M������ҹA{�d?��eU㘔�=5FށՊ�`^�-C5���Z�L6E�{���0��Rը��W�g�Zҿ��T(�+�<'#��W�IW�h�9Iy�؋S?�RL��<�Wo]>N����if�8�䕤����&��i̔~-�J~8��������y�3/�F29��6�1nDbFԝ�����W�:�Y��ƛ�	��	m���+s�~o�u�T���;Q;�2�C�k��*Aj����P<��+,X��{�/g��������`x��\7��D�'D��vr{	m%�\6��V�q~&ch%@<lݏ���Q'��93 �q8r��8S�;�Y	��.9�=�&�4� �n�íَ�8#��i�U�6aD��'h��ɻÌ����2��v���i��V�L3��:-���s��o�Xyk��+�0���X��ރԃEσ�Z�$��~��]	+�\ݦ�Ro���t�.oI����w)Xzz;��sg�=���})��~�-���c�G,^e���:���(�C�z8�����:(����Au#]���uY�\����B�����J��^��(&����ݿ���Ր�YޜrC���;>�<5�fξ����$�'����vNqcU0ض�m;���:�B����؅�(�����Pr�wt��z3�$s�����[C��r�w��?�~� l�N�51�.�,���ȕi�^4M:�2�Os�*�z��5��C�6O@tPv��)����pu[@}���E�#�U*�̟����ft��� ���$��% �k�ߑ캁������3�{$m��m`�D�HGU�G	4�\�l0�ߟ�i(��gl(�Q���N����3���H���%����}^��yx�#��跾��ކ-  �
�F��Ѿ ӕ���	iy��=%
��8{fe�\C���6�*���EuBq�׫k{�A�`&R�z���ΈC��)fpQ�L��?����7��XU8������{�9����%�LT��#��Jz���Ɛ�^��H����M��f��ϛ��csw�z�4����jjB��Ȋ8�39˘�ճ@�rĎӮM������j��ܪ�(
�"��$9����ݚ�#/E(�i���ق���w0iF��V1� �(�N��i�9���4^��g:A� Vg�5<�(�h�/\��k|EV���=���q�tqk
�G��V��7|����S�0�g}�0�(�x:�5ς�_t|QM*@�/��� x�E?����C�tZ3~#  �?-�-���B	��{Z�)	�v�}C�AoS)d��j�Hě��4�C5�7۫q�DŵB�ɤ�����LeH�6W+���9��'���t�갞{]�L̃j{j�pב�+I��_���Ɠ*�U4j���+�bKj�w���>I�V�Mf��U��dN��ū�Y�}��BB�=,���	�kߨ�*1��tI	�#���P��)�z�֣C�+D}ۇ�>S��G�&�b�W�:���Ԃ�u��7ux�������}$�����k���&�����D�5	/�NH ���_kD(�(�*�8�_�}���ad�X�<7p���o@;mQ�P�ލ�����x�k���(`�Z3�#ֲ�@�ΰ�f蒈v��GH�b۾�l.{�JR�����PE$`�� h������Zq�q8pd��]�Ç����Qh�(��dc�LT���ьYprK��iM�X�}e���� �k=�Q@a�"C��S�˥s�ߎ���ΛpsAL�4����C���t�)qc���t+�7h�Lcm���wX�b��B�5?&4����ku�|zU�%[��${����'�y�l�~�ζ��8�k�S2V5��e]�:&į$]�O��R0���N�Qg2������/P~>(Zn<�}1�I�����v�13�ϋ�]W�9�O����&⹈�� �D�v�1a�Pc�����
�v[F���ZS=j�����jW8H��Y�a�D�0�-T�? ȹo!R�{f7Y�*������as���G]�8�Q@T
��'Ww-R�����fP��9�;����>�~mG*���3�����ï�&�l�T0��b��**�y^���6�ۑ���̒y�O��f���������>œ�t{��zS5�/�HpjKk+ƅ��+o�G���[kR�j��}�Œ& F�����F ��^�4��� m�^�"�4 lد�P)$;�DD���?nk��V���sW�$��	����nа���|�3�h�\d,c\�E�@��������o��}+��=*r�f����_:�Tܟ��<���$�w��)Pc�n,�p3e����?�t�3������i㥩��w�m�@�;g����3�僽ˇO������>�?�Ȭ��}3�rbӓ��D΋�X/
���o�����@�����L�ܬ�L?7��Q�_?��R5kÿ��+����O��D��#����sŢ����\���_�J��+D��'�d��㔜$$��ȸ��=��#�R����z�;ۆE~�������t��;^@3��-//�a�N�`F��_�3{_���םeִx6��$��XG읭sӻ�MdB�)9�Y�Խ��$�kZ%)��d����P����R_�O)zB��*ӏRŭ��w*cEת�ɝ�|5�<G���!�!�tV�(�u{(˷�hd�1Ơy�^��Tæi������3<�N��>V��k���QϠ#mx�O�ܴ?������@�l=N!��j�I>=�FgF=���L9v��4�y��?�m-0�Fi0��!��vz�I�CNݺ/[�F�YHϮ����zw�umk6Ts]�7�_=�X�m�(��Ld{X�h�8����+/�Ww�9M���4���� n��&����8��9�E���"�����Oi�^��
�R��e
c�����}�ddT6�I>���z~�%aBZq�r���SIӋbG�Nzfe�n��b�n �Q�T6��^[�d��L�T\���?Q%1>9�� b��,�]`���Ilå��OD�0!�[��W�ԵE��;���ө|��].0F+^�GjN��r
yw����;K���~ˮ̤�	���y�Y�;�����hqI%�i����d�ZAo�@0Ǹ괄�W[�b�T�?I���xcǵ�X���Z��O�)S+�}[l�rlC�`��������k��b��G`l�#�<�Z�5�mE��d������[UQ3s���'��rPB���[��ӵZ�
b���R9��x��K%.C��~�ἓ+��TyR�ݯYU����f�^\Ѡ�&\9�*�j�9Ib���擇�o�t��.fb�Wҍ4k�i_��m/�~�'��_}�H��c9ؔ�������5N �a���޽{_�R=	S��� p�)�$�J2�/P��G��k6j-���ҝ6��.V��K��QV��A|�*��<�r�M�3���ͱS=t�KR����?f�#���'�]�v���Ic� Orpt��z���9�ǇYC�n6�����7���ӫ��T=����D�w�湄��q�ΥM/�h`/�Ġ;���u��"��[��Ņ�0n*�C�[7��_r��c��U�̪]i�#��b��X����X/��s��oז!�L"�b�8���ݚR��`R��U�w���t����1���� � \����#�?���#t���|��DFl��t���|��� �3ؚ)�c������'�^���r~I���:�Ffi-A?��g;����۱�����е��3��Ӎ,j��X��^�F�#ݣ��^�,tC�2�'~���Z�$'"�k��]D;�z��r��`�z�.��3�!*�Q�R�ҪY��b�Jbq�3}`T��W��Z��"T2.\=Y�����ǉj�{�G�����N6}�y��	ɡ����$�K�|}x܋lr��Z&%&�E
�kٽ/�X�u'V:�Ø���I��j�<s%��^��G�:뚤�6{\|{�QxJ���T�w
t�*��{0���Dr��Ӂ�{��ڞ��6_�19�!��+�5��2cV;1s����/��o������$�(�[#�u95����u���0����x]��8	'�y��� \����U<�O`6O��a�z���ʪVP��B<	����U����Gh��ABڥ� 7FL �.*���;�f6��5�4�I
�#_�S
<��c���K���1�Tg�	i�tR����p�칤��`3�����ɯ_K����3�=�w'��R�Fk�O.���Л�e}� J�/z۰i��crX�=����F`M��1��5W�
������91�x����b1�&��nK�3�eR4
��ӳ�q��p�����Z�Z�lg��&L��F��l�Ǆ�z��5����MZ�$��u`�G�Ev�-��+1��s�޷�=o�/S?����p���OW���(ibYf��n���xv"
^�~�6x�,V�=:;ǻx�87�=��n��V���dne��ɠ%����(]꧐���G}|x�v]�܊[�@t�� �E��G�l�Cm�6l�\�ӌ
㯝��߲b��
�$���Q�����r�z..ˍ3�R����H�ZL$;�rs���WDQ���j<��Qα{��vD���f䮩��$�.�D����\gK���ǣ^;�׼�a?���:��ed���*�%�������(&Rt�+������z���O�yx�\t��S[�GS�����#w���F�O}��݊�J7�%����X{�3ǒ�a���<�cS���3?�GO��y&��	�
�z�v.V��a�z$4j����$�	V����Q��Z���\quFG�٢��w�]L�D� �����y��e3�lv�# @ƧY9��2��2i��z�ğ��Vn��+	c3"NO�5G�w]�V��E(k�m�r��P�O��A@Г��!�,�Ϗ�S�b�=P���(d��f|c�K|��t�^.kވ]��cK[���1��ݽx'�.+�a-������$e�fxӿ�����B]�T��b�u�-���y�Y���3/6�86�?���?Q�FY���3�M��N���<d����п�T�����Oܝ)Ȧ�%�{v�l>����q�$����\���(\�Ys8V��� �D��Lr�M�Ȼ�:ϭ��z4����qh�دy��~-QT%:z�-�MZ�@-������,�*7��nzЈIarR8���K�2,++!:�܀�CeE+�?کI,ns����\F��Py�o�۵@X_����%p�(�p��N��qb�Z^m|��Ϩ�B��J��'p�P�ɪ묥���ׂ2TnH��u��t4Km͌��R�+p�����Կ?��7_Uݓ��	{�J�&m�W��K�{�c�$�
`H_d*��0�s�x�%#`GeMp���b�ʅ������+3�|�\�O��"�r�%#�����bx6�"d��p
�ar�[������==O�>���Y��1@W�O�ԛ�&�K�|����Բ�>v��	���������ݨ�פr�ܙή������ǋ�]��	q/�_��Ɏ���7,��!������z9؅L��'��;0��ZĹ�-T sw�]�}=���b��{�k�é�xm�v3ͭ7Q|��,���^�_�{/�=:|��� j'���*��=W��d�꽥+�+%^
>�͔��a�b����}�ۡ�ҵ����"&�������Ŏj��0�ˍ��J^r�O�;�pE� ���Տ�N�w���U�S�gp�)��ϐ.���4d��Q����s��]CÅ=�O>kF>������ڨ�'O���3�bN�ѵ �v¥�~�j�����(���ӫWߎ%ޚ���8�9qlz�!4�3��y�ɉ�Am�K�ԛ�}�\t�\e��Y^u��#����O�!y��/}���Fʬo6�����h#�M���;�\R9,�����E�����;fM!�u���o���J<�]����1Q+)�x��AB��?^�����!DF�Q���s)j����o#agZ⡙��*L�8C��a�H�3,�@o��~O@t~@u�jW���U�����-�����	T�7#}]�EY�h��;Q�.-�~�h�۸���/!����SPK�̨����F��u^�҅&U����r��Hr(ܕ����f�`�s�@7���3|�t�����
���/��\�do���ٕ��1��.,�1��7�������Q �egU�P��ʒ��Q�S�L_�<����M�%�F���%z�q���9����o͸�؇�h�uy��
9�>,��Hw,��S��8�δ~x�����Z��'R�1�Y���c���l�S��C�i�C|K��p!�t#�ߒ�2�U���/�4���ߗ�ie�1�����:��S�.�^�or��EW-��~�sM3���:��t����v�G#��74/��jݙ5�ҕ���C���"#���|[��Rv�M������Lu �f&�
	�d���g�eR��t�An�b���un���Jz����&����=���t�tYy���sB��Z�II�\",�����c.���&չT2
�y�OO�Nm��aBX��q_�<��G�yx��
:�Ȟ7�J�ܸl������&Mɍ�C��|�XNx��#r�+=�&�9�����RS(_�.]u�D��N��4�"����#ل�:��΁��kt��V
9I��P��n+��7Cr{r���o_��{k�M��w_�@K3z��;܉�J1�o�p��{���(+v���_~n)�h����$��p�Wc>�}�d�oN�%�]������4���S>0�H�D�-�jל�[�x��"�CaN	�q����'��9g����<�֖���p�P��ZAQ���U�i���9���XE��J�+��&z�H�E�����w� V�+T��dϖ����Nl������&n���_��W�A�	�?!5"�г�`L�)>�y5|5��g��-@����kj.���V��0���� (��\���5��7��w9��n'�,���0ڧ���(B_ �|����I��۱��s��w���)>B�}�ZtK�`�_��ʬ��6����2����2�J.,?6?/#�؞��>��ݚ�\5 md-��ߢč* �@�M�.r�C����`���XY�(����s��-�9}����=�A[��6��0����QL�3��b�o�3�(��_��"�:dJ٨��n^�$�?��!cPW����D-=���,�q8��VN�	�/Gľ,��\c4��������N��uN��m�؈��d�dn���M,���b�m8�w.��Kg�1�Ƿ�������;�{���b���_�������L�R?Ңv�C&�I?yK�9�T��|/'}ǽw��ߐ��13��u7�>u�d�Q�=��7M��h��-����jߎISk�I
6l�Z�����Aᄾ7Ws�!�뒎�p͸��$��\޾`��>��_n��>eU���	,�ѨTB(��J�9�v�L]���0�r4׳Ԅ�S�WiE2ڼg�#�w��PY�K��l���gZ�=-M���3��E�7��c����n�)
��IʵJ�7�Q]{p*ft�삧�'��$& ��R����q��Pm��Dʛ�>�/@���&@�,Y��J�,�V�~����R��,YH=]O���R�bҌ|9�['�lߎ��z+^����zq<%��Z*���zO`�mߗ�6��G;�l�-�ƿoO\��Ν���~�@�o�J4�h��	��*	_��7{�ydvᙉ(�H�f8��zz�,�����)�h+*����D(�}|�O= ���_�xԉK��^�m��oz���f �Z\i{�M\��x�
�"���$� ~�m$�ǟ�=R�������֦�����N�����˜�Ǫ31I���3����k�W �>a�(�ܯ��4���no�|���� ��A����J���@����8�窿��T��*5�0�k�5�닓��^?�+s�1�%Tjazn�`:�C�Kf�O9z�I��*�?�R����?W�+.]�ˍ���D��w���P�'kL��w�2����]Ւ��%��R}���.o����}0|��*'�P��*�0�y��g��WY'��9)?.�����5�'y�יm܏KG�t��vyy9�mV����&�[o�0@�r|ޏ��^��V�E_����'zBW�]Gt_�w��Hްi<%s�S���6S̹�8�3��l�����;o�B}�7���l˵��{�M�gXZ,����{H�[�)�[V���@�cip�9���7����1�[�)�����h�{s�kK]eO���˽��^�t��Rz���\�A�E�nQ%������ɣ��$|��QS�_�r���r����:�ݭ�Cȫ�7�������g�P���
��rZ�33�bxT���iӶ�����
QW���;$�������q���DI�&8�o�n鉡F�ς�j1-���Z� ��7ţ�:9I�JL\���q�*x��-Q5�H ����{�ܘ��%b��_���DJ�SO]�jd�5���0DKw8��Y�e�!��fиDD�r�,�Da���Fԅ�/����Zr����z�.���]_��I��o�xS����¼2�F,�~9i���b�4E���V�gv�X�a�I�אJ�C��wi�m[��vJؼ��	��x,Ǥ�^��A�/�6)�^�u:�ű|AB����n���iӠ1�Xa�k����a��.�fNqF�o��^��?Sn���
��\n�%�܈C�@�fp8�� �V�8���m�l�� _(HH�H��R�Ҥ�WJgmm-�2`�����>jz��v��o:���_��k�~ʺw훽��gH���|�.����AR}fX�,�,�7PS|�p�@�Y�x��}��ē] �\�V]/!��xD�˒&���@�8	Ԁ��_sݳ�cv��f3S���[;�$�����^!�h���4\�78�����\0π�XO�����i����KR����8��脗̰�È#��<=٧����N7�̾^ ���Dp� ��p�b��� �^���V�������j�v������o��ԙR��J'��{>3���suU�tM#5�I�̹ܿ�o#6��f���f�[Z[g�+�� ���H�9���z��.A[>r?������v�Tb)a�K��:�`"j���I=��"&^�Q=�y�V��++'�t<��+��u�)�\X�qf��Es:�Y�q�{b��L4�n���F�'�h�� �$)�|�i˙�3����$�*8��/	�m��������Z���ɇ?��c��q�\�����;�S�G�C���5T�u��`b�i���h�m���5�peŝ=���[������Y/QDho������fg�Ż�j���	ِzj�N� �~�]�j-�`V��$���
�پU�o(�꟨��V�2����cjm�{���D���;E$�(��˰_�#<�%%���@�`0eeev�b��	�
>oQB���Q(4��A�(-�u�� ��H�����uuu7��	�9��IRsuuQ�J�7;=���k�����vƑ
�s�kc��v��F�d�(�3@ټ�_��0O݃*��=.��cg-NA��G��,M�n?[>�XNH��et�drF�Q���ٸ)��M*��D���6�㰬��� ��W��VOR���~I;V��r���,�8� �'�ڰ���~�Y��ol��Lg����q�
;FA�ON	8^��*�C��~�#�镍>����ůu5�\{d�-��s���p�tG�Z$�1���3�{�Ω?7�u����f�E�;+�|��9o��_��KikS5m�a�
&�Ծ�Ӱ�u���#��5e���D6i�V)Q��K������z]ԇy�@K_���O}�:A�pz�
[����~v�Ѽ�����$'K�kF��4Ң�%�S��8�h�$靯�dq�xC�7 ��o��8�т�Ƭ"��n�D�93 �u(�t���d��ʓ�T�n�{�o�震ө�������I��Jt���8�6��|@O�q�q���
����/A}����а�cN��{�m���C@qH+�h5���U�Ͻ�mQ��ge��P�햣�a�ޙO�i���:�[�S�����=F� խʔ���~9��+�}����i�6�q=�:C���-�NϬ̤�H�Kz~�AZI��s�tҳ�X`,�p���u�l���u��:�J.w�k�{?� Yz* $���"U��?�H�l+tȼ�{I/^�H�.���|�=bT��ՄrtC#åay�������n*J������1x	CzL�c���)����~: ��CK~1��fxb- Z�P6[�VPO/1!a"V���2��&5	�[���ttQ�(����ʏ�"���[չ�<ak��)'�/7#��:/*�ՋO�;�J��{k,%���_��;��&���C�7:w:,ײ��,y]tz���;.䳸��w���}���-�!�͞�Ul^?O��C]ɽٵ� 䱄n��D9���)Ig�SĜ�ڦQ�ib�K���o4�d���j:���>����C��`���Sϓ[ZZ�T�x�@���'V�����J(�I�k���)Q�S"�����p��ɒW��b��������)p.,!���u5q���W[lǤ�Z�ѕ7�*��T��J���ͭ����!��ŉ�y���|����*��,�]�y��UR���� N��i��z��r�	��d�k)�l�v�	�RYr<)����#7�����>�Bc|�V�B(<0�M�����5���~G�d�@�%�h�6	Z4��p=��M��ߣX���9i"K�%�ENm���eH�O����I�n�zí�Ǐ$�]�����J�e����_��,���94�H~��.B���k�[�D2-ׄ��8 �j!�o���$0t������~�[S,D����m�zo%)ʚ����ܝ�}��[3��n��骷ز���@#i�Yt��E7�+���~\\<��u~�f<{]����Qp~���V��zw���P�+P�\��(//?�����d)����-�, ����,��\]��c�1uBg��}SO�'�����hF��P<˛!��3�S�Ų�O��qBt�O�*}����̜&�$Q�&�Ukx��j�ʹ/7��';���w�Eꊥ � ���L��0[(4a��/���Dmꔋ�>��_OZ�)�$P��ꤔ��0�¿Y�8�d���������Z�o,_	W�U����M�y 	�FH@p�$Xw�m5׿4
��Y�YKK	sZ��5B+���&Jm��q� ����J5�C���2^ũs�?��.�Z�.������YU*���9^��
>�8b�:[v�x,�\a�|�1��p�������w�x	�_���=a���2x�m/ϓ���І�N����{�:�z~�B�7��ݑ���?%�À+�[��L��ܻw��֐�<�����r��W_���+��G;*�R�`.�9�mN�w��vأN0��/d���i8 ��H)շ��6�/����j?�*s�����)�?�o��!�b���a�ˤ�.��bM��m5�������%���s�p����T�r`�i|�3�l�}���u����S��W+-3�=��tN<<��������Ԕ���Y8��A�Kg�(8�v`��X��87s=ͷ���TJ��,p�t!�ك_��F��������ҭ����ߟ�����U�g��7{*��|���=��d�R��hH[��������?#䓓|�sx����f7����Pi $��or̿~C��F���v4�F��chƄ��HK2��viS<���y��g)$�f��7CqU����\2Ђ�ŰN�k�`��\I<��%E����v9��G�ׯJ��|�ه^y.��d���n�$ ��ں~kI���R|��G�x�����
x01�F�b؟�%��?;����?WW�S
ǘ
��?U+��3�������	���/(E�ė��~�:����S�j�P8tB��VKT��`u�k����R	�%��a���� 礊�N{�	�Z1��ᖑ(j�o8�OvV�+��P����U���Dg-^�����ƺ�uW5D� ��O�kmXv=����ǚ��-m�ʪX��f7=S�jz��L�K�dy�����B���U�mArS �YY@����Llm+�GX������s��^V�؋�>&R�5ꏥ�h����� z{�PU�q�a刽�C���;������߹5��_�U6��c�Hh鉡0�Y�8��N��6Ѡk�.d�/M����R��J�B�q�׶�������&��($|�g����y`_5+N�ț�s�2����2�e�=t=z^4O����bB��lwtuu�;��~�`~_�S|Ҟ0�*�a$�gi���鸤t�U�q��.S�9Z�{6�,�������'�?���9��%B��q}\r��ddO�V#�E��� J��A������{� ��p�铄 �9�k^g�LD�����jGzI��^���ʀ&6�[�����=~�ީ�
��W�W��SB��g�e�qfR��G��Ȟ����YՇ���UAqG�	q����T*i�<:x��r�0�@`�Ra�Kg�_NV��)\��j�����<]m�y�:�N��S�M�|�A����ĭ,��t2L;%�p�q�=��``
�xJ�9䜒̅ݙFҍ��W�t�z=�|tA���|�K����Il�'Lm�)���ϸ�F�0�|�.�{*�_D��b�t,���Q��c�B��_r4p:|;	F�$�ܬ��I����M�az���Us= ��"I�ܺ����K�����.�.�Θ����(�F5�����F|�_XE�!���� Bj��Й@AdS֐MЇ�(k�Q@��D���S�߷����%�ˁ6+Hg\��q�g�9S\�s`	��<^�")"XE�^,Y�<�q�Z��.p�=�ř�fg-m�$x`�٩�~�( ���љ���L�5M^���49��yP�=U��Ȃ�{���>�'�F�9�L�r{��P9�i�v��S��\��[��i�R�/�Z+�xGP��[�K��,j`��������ݚ�Z�V�Or�K5�}���]�*��<�O`F��f&��`���M_[d�C	~���J�/�H޾~�^=c�#�-�ܶ��Ҽ��,��9O����<F]���2)�4�J��֜"����ӵ=��-ǲ�]%Is�����H�ӎ�;Ȱ
'3�+N뗨iiQ鴾������q�X��A�YY�LMO�l6����ZCHo­���(A��w�,������F�c�>���y���e�5v���ֽ�^�����
�g0��{�`v�#D䏏�\k�^Z���v{��Aԗ���x&w��|�_�\�;��f��.�k������/�4h�3�^F(�$��3�FA���!��f�$�O}�/�Zd�b%�0n��M������p�ں:E.m)�z����30@y�P�)�RN���2����Vx�_��أ����SNQ��7���q�.�����=�Y�ev�\�oTR1�'��F}��Bd�7	��xĻ�*׼	�{��=Nv����z���k�������e����5��(�;u����K�(B�
%2�,Ƨ�i���'��	k��<AFH�Zwc���'/X�i��@$kh�������~xI���2��%���'��/j(>��)�.+/
h��2�Ww�0L`�d��K�W���Kg7K�kF���O��q<Q�*�w�6)D�k����Eo{��A��u\�>~���%|M6�@�"��R��[gVsk���T�����ܲuq$\~t@�
e|�3�m�6e$���WO�&��Oᣅ�kr���u{$G�p�����۴1��14"�4�K︌kt�VWl/��R���L�F_aǜ4�Uq%�U�����kC�����+�>F�~v��镉S'QWD$�9_f�Q����t��_B_��5�s��� ��q7S���hW���^��hdn0{g�.���Q1t���hIq�� ��	
)��l�H���������y�{��N�T}y<����R���d)KHc	�X�o2v��:3��,�Ȗ%R(��ml�m4�"�5�$R��;���|��_x�<�r�gι���uݏ&V�!9�l�/P�j�(�@ ,��-���?��:'��ߢ�7���:({�e'����k���۳1u�͙҂�R�^+J6{� ��V����s�k�1\z��=~�A������c7�����E<�$��Ũ%grr]��!����lҁ_t�D����2Tm�� Ut�^�4�X����ݘǤ�]B=���~�jk��`��Q��dx�F �: $�yf���Z��n�45)���W��>4�#�XSyMY��O��+K�A<�{�zdm&�����e@� y����0�ˮ�=pAO�nQRb��!�}����D��Ȭ|��n��,�X�n����U-U�FZ\�%6vvy��r����¥�c>5��>^��!���3�@���������v��X����V�3d7�H���2C������G�9��UK튤���x?g�}|�1hz+o����(s����L?������2щ
ꙥ��>8Xݒ���U����}q������z��0�_���l�>ܚr.���X��=���JɅ$���;�!�I'dW�ѱn�M߭��{�W���Vp}�cNѹ�2l}�N�΃���͜Q�^�	�=�{��r�g�z�k�����j���Iw��	�N�������:Yw2@�^�M!�=�l��`�t����)�����b�ș����)��caU����l* �{t�~��I賕Ҙ1o1�/&"�UUG��tu�ė�����'r���8=�~ ��|d�~wW^&K��Y�D�]�1Q��1E�*�)�� �Ѽ���V�?Ӡ�W{nk�ȗ�&=�K#2��j���]���|)�,U�C�r����!9���0�y��r�]��$�(^c�Y`�0��7��-3o�K��bn���o���7�o1�4o�Ɯ�L����l��zyl��������W\x7B�d˟�:n!�e���@;�0�و�T)��zh�ё�헣7eVRЬ�b���W�����ͪ��ȏ��J�����Sp���4��ND���cz��y���� JĢ�SW +Ұ"�VD����>�"��T�y֪��g���J8c�`f��B�ףt����KB�Y�)z}-T�M�6���_�����%��>��(뛇3���ʛ����P�SoSP�<������R,-EzG#�ݻ��1��[��1e
��	��Rf ������K� ��n2%��@Uh�m�_ �-�؀�K]���Q{���xz�xL�г�� �Y���.~C��i��؄�6�O'��5鿛^�,�Mg�{[u�����Ϙ�1o����ܯt����a�f,����1�t�3�8	m�P����.��|
��#
�go�����+$���5׃g3'��g~G|߱��c�%�"����j��ʀ��S�L����L���A��"�����ࣣ�3.���{��=���%�	
��9$��Y�^�}�+=,���ڍV�?w�]�h�s,�%� ^=:��!���+Wk�4|��Y P��<���"m��Of`��>��ϭ��F�#�����#)�z�usr�HfT<�F�R��W<�1��뚬l:��T���x�怗�J���S�W�}��"9U�o�?�f6^��0��!RG�G���$Q;R��}�r�<��|�Q5r�]Pe#DH�G9{�O�)4��,���s���A	�u��D�O1R	���O"O�X�J�T���d���w
��0g�7���n����ӺX��g�w����|�A�`�t�ܪ���od����6�������.���g'	*H�/a������UL�ߝ4SH��kҠ&�
�$���^��v�Ì��e��ǖ��_�#5�ݙ5��_��.��`����θ{W ���4�(٧�L��ViE�th�����_���� }'��S��wS��9a���������������cY̿��I�2��El~ܩ��g:�"ى*1�\t�:zT��K�ɠ�����ހ���6����9��;�d���e/��5݀�rj�eu!w@:\9���tњ������շs�_Y����24;�����6z�Q�k���>68h�Ȼ��ƨ-,�#~D�{���ϺP����)0��N	7���Lqe���+jrr�:!|g�|��;#��j/Z�$zI�u���Sd�Gd\�an�&�/
�m�|�`Q<x��瘸M�ٝ 3m���lNFV1�N��n��R�S��Ɛ>_0C� *�NQ��J.�H��J-n)��x�B7]�4���[�O�t���#Bs tOɁD���xIS��&vO���;V��-ώqE��YL}�
�U����(:�<;��O%wa���G�	�lAU���x�ɳ��U,�C��d���i����%�5qQ��>H&ѣ��0H�W�����::H�⩆���pGK\�
^���G-g|.���5�]�`��lUK�p޿ױ�m��p�U�_޿�mow+�ͬ��3C���������T�+���b�c�(<��sC�}<���CQx��އ�c�1?�d�(!�nR.���Ŧ�\���&��i��&M�\����,ӎ��M�2+�T�����}��n`��ؒ~��*����
���c*�#)�չ2�1)�$z�����p:��3F)8�Q >]��2�皛���@�A�9�A���Ìd׈B�>c�c~Ӭ�ev�������ֻ������iт���Rl�;.]�Sz@5�s>�h��A��C���O\8�])Ma�"�	Ji�ů_��uB�LMNF�`z��i�M�����`���v��Yw����h�σ�̰R:�-	��z��\�2_-0��W 5L%/JsG��AQT#��>��Ǽ��)?r3�9�䝐����z���?e���h�/ d�wJ1b)�׏��҄���5=A&rrB&F��;y�U�c��\<�>���WO���-~ԙ�y��v �o�V�� �ŝ�4��>:��D�/8׏0��T�(�<�D	��V��B.���sun��8b>������E'�����E&}�>%�6ؕd� ��\^�Ǯj=5O�����=A��&�P�D{�;����I���)�Wv��� E��sݾ�L2��]s���T��#QA�w@����~Ij...��ښj�?~�<���'T��K��/������ c������x|�7������^^��rqV=�>�f�v��-�s�yJ��ߖa_�(/�4�����ky����]x�����K��W� ���?AX�vab���ˋ�j�LZ�6���"�וkL4�=D$H���+��ͱKxN��	�|d��(�p墻�o�)�vY��ZyC�_�N�<41_;�?Rx?��8�Ae���O�K���i�w���:��P�$c����5́��4[O�3�^�v�¨-FT���:�/�|��-]�q*�n@���?�S��7� ���xYm��!��9�W��m��&�w�x�ѝ��)}0"8y%k�����9��#x�<Kcqj]��Uu��۱�ýi�m�d�Ӟ?��l)�����	�&j�RN*%vܵu�~e�ߢx�=��=0��ۅ"mY	���7�]x��>$�0���^(}u�Fz��E�F��G_��b�<�%]�EF��|W�v�#0H�d�ŜhL���s�m
�ԓ4����H������@���pj��3�q��he}�,O��P[¹3�J�Ji-���B��[��6:sҏiWv9T���e�H����)�����hr��w%S0�a�퐿��䴪�y�d�p8�IxIb���J��f�92�ܠ^d���~$:�O5�itQ�i��~.?8�a$�V�9 U+x,}Iͭ�̆���<�f�>*�V�1���.�m��y<�f��K�����M�^m���'ʗ��e.Wu���[��\�ߕ��S��XK]h^���<F�Ң�^J�/i`�Օ�J9kACTT��2���R��|	L��M��idDO��H��VCcl���)dX�I6|:`�Y��x����x��Lcpu�MےL�at����gMVm���R�ג��u�F0�k�j׸��>��} � �@f�&2V�a���E��GD���8�T����`�Z�}��'9��� ���U�)ck@�s�:��͇{����ȅ�ia��@� ���-��(4	����q�����2��V��W�{�����b���{BAJR�I��#�=,w���s�[��2������E��z�6}��$یd�=��a��V�k=������~vm�_�>	6�țp�tx��=�Q��؛qg�I�]@bջ�������n���փ�(�E^͕�������LV�|,M)�4���r�92�C�!������"mCG��Y�[�){�)�.�2����b9��!����� ��t۰�j Q-��޾;���{+���M"������P놛,��jp�\�����/���N|.i�fȅ���O1��O����t��bo��p@�USW��3|�;'Uģ�����PΩd��cg����L�d�woa�u��$�'��k�b�
��;
G3 IU�W	9�m*Pm��YJ��Q�XH	5����\f�������A���"R�j�#������o��-�#k�EԌ-iK�߄����ܮU�t���},N'�ٳ��܂��B�@c�j�S$��٥���[c��@��1\"Y֭^|;�r�C2�9�3o%r:�q�C��Gq�/�JܞWIU�� l�S�]�yv�o�#E��"&]�?㷁	qY?�q�Q4W�J�qŷ�x��Z7?�x�'[�	�%�c����tF��R��N�����f>�N+�M��N;�;5�n' ��r��7/���EJĝ/]�߲Cpl���|T���:���^��(0�"�2��C[;�t�^���\���yn�,�󗘝Ǘ]>C�pz/��tr���	T'�������b�T!�\L�yzI}	�9~��c=<��k���5v��JF�9(����+>7���Mk壣���q��O
�H��FGES	aÜ���e���&kI&�"@�= �X�"e�)3���򗹅?��D� 0�?D��:���ʨ�J��H�t�������tb
1�1�bk����<���&�L>�v��=�@1����X�I�Ն�_��۝獫�E#8&˗T�{'��A��?{m�{�k�l��5M����;K��sh�U��9<C7Y�iz�����䭭�����{��pD��������M�<˔���W�3QY�T�1WI�y���r]8�'�0���).�B��SM�%�JY�E��?'������-��>�y�K����R���!V=��a1�C���)�[dhp5I��k�z�PcC����k�:�/��y�2'�T��Y�O��9��ԺY[�N�����"�j=�|@�	�V�g~�E��5�O��^��Z��Yt��)L���Hȴ����$����x����]��\T�Ǝ-ѧ��%]�2���,_ꘚʹ���s��Z�Ai��nX�t�~?,�������=${��^���L&3x���0N��	����:n1�<�����~	"�N�6�
�n���V��2�4Zԃ��m��`��R=�r���X�%�_p�y�&�
��"b�}���'� ��Sb��@'p�!��̲#���4������w����s�~\�?���(�������u��;zu�ꛊc���<*Ty���)R0	%��â�w���s@��t�� �V�A��t	F�/��ۂw<��F�m7����E3��ջ��^��� �^�h��ꃚ�M+����=��şt�JA)���G��`��J�v��Y�Bz�Y���"��|j��'�A\Wڻ���Y�%l�C���տ%���i�R�T�?��JB=��Gq� ��� 6&xEN�c4���m��������ѤT����#�>�����=w��]'W���JL|1�1���@>�^=����Q9������`�X�Q:7�9�D�c0��xg�Ջ���"�y��k���7��!?�Ћ��X⳸w*�8#*Xz� �b���t�/1GD\؇s�q3Dn}n8NG~z+=L�;��_!���������D	''!�*�{��[Y�[�j������l�L0�~{��;���YQ��Nz����9��n:��/0�*
%}x�>������`sWܞ����({>`�)h啰���"+G�O8dę�X����|�^D���y>�iɏ�r��S���P~J� ��(���Xw�h�������M���I�;6'���O��]���P���Z<�Jm�:�,�y��t��alb��9�rD����=d�-c(� ��2��3�H��
 M��ySJ�b�;".a��P�ቀ������قq��z�-�E�I�r�A�I�^H}f����f^�&j��~K�u��R��|6���sُ
�4�����2�?G ��ypaY�r����}}����h�s�?5b ��?��M�ܭ"�(�t1�[^����/9�o	b�\�'�,���Tc&˃Ԧ�}s���!A{K�7l}'���0��TV�z�Pq�"%\��َ���~ђ:�%
(��g�*��㦽7�5�Ɇ!������Z��Ů��[��Gd����<��ԯ,�9U�⬁�ֹ��wݐ�k�?��?���0�p�ZnM���=�w��9� � `ޥ����ru<_�ŉ>b��}#��s'>X��PT�_����]�V=��76�>��H��tr���<���}��Rl{�8t���P/��!���/_p���j���ܲe㑫O�L&w��d�~0�o�$#�YA���{mӹ��|�6��~ޫU��!��)�����ME���Y&�
'h{�m:��T�����4-��?���Ǻ7f��	��UF���^�\7n��g�6�ȯ����"!?�	Kټ���v����--e�Լm9��W��Aj�&����Cj���Q~�._��3�S2.F���B�A��@Y�WWWuO��p��U��\����'�r����q[��u�\�y��D�}�wGpNo�2��viga[���c޳��]sW�<���#|a��ˮI��a���C�����)n�]�K�yk"�td�].�myֿ��w�!b�0#P����ׯ��^�x����mM���-y��T�_�ۺA�I�;�q<L4����[�E����#ù5�@𩐽�hf7^�������^?�LRg��yyjy��� I�{*C���^��_�?ǡK�6~����<^�+� �����-��Q���>Ai󬻻{���?�^p�>?A�a%�� �����qҰ�f��H0�EH��-I��G��Ə&�n�]p�6�B���ݒ����'P��Hq���-������ܞ���o��M�����a�7�wG�ߥ^���4ܸ[T�7�E�e:��)
�n���	�B�"K� \��ZZV�~��g� i
`;��C޺k�OvRh���-��ɬ�9��A�C_��E��������U�-��j�;�J����	޹�T��� �1��?C��ِZǰ/�
�S��r��Ĩ��fؕ�A�y��B衭���iҼ	.4
խ�sZ����uJ�M�$���M�C��mk#�����z���8-K�c�(�_.0j���$@�k!�S�i!�ID�C�TQz����-}���AD��뜀�	u�/�ݛ!?>]�������� ���1�?�7�3�NÛF�X ��3�\߭�騞����g\ذ=��M��෉d���@����O�p�S�_c*�D ���k�J%����Fa5-*���	�2���y�/��<���]���`����w�N8o+״?j�U0���c�J����0�{c�L�[״���~!�M�X�s���������P�ftil��w��3���v�����%� "7�HBiM$�#��U�Y�̥�SPr�1��OR�?m��蹡��2s���(.ew�m�珀�g��:�I�"�����K�>ӿY��~혓��96���+�����w5]>ɧ�
l,Ӯ� @���p`6�����e��y�-�"��Õ�S�)�U3�It1d:Ư�)Q5OҺ2�c͏d�� ?άh�� �?K:�{�GD��~\�����<X���4�W�V���mzr,٠�x��9s��po��x,����Y�(��ۭ,\\\_����(�S,��W��TzuF�J5^�:���R�q�B���lZ��5���-٫QP�Q%�V����\Z�-�/�x�?$��Ĉ�1M�y}c{.A�ņ%����VY\��Sr%�5��ap�/�����Q������7�J��}�A�B�%����f\$��2є;�X���1?פg9wfO�2�~y����J��u$$���D�qѱ23]����iI�TH����WGXN�����ٳ�8�J��3o?M�_~��Re~�����_�8/0P'\���NOZi�����~���ÚCӞ�9���̕K�w��n~M��Ir��ks�J����vD��DU?�PJ�}��rr��oC?n���d{��\WWWG��˨�/����L{��?�5j�t,�I6��t�M�G�u��c�� a�qb�^"���Z瀏VU��O��7�u�}z�9Ϋ���ڲ���5�2�USݸNRVZ��ę�)v�}���-��\V��~�1�@��J�����m+MC z~}w(�!�z�A�dΎcAi���4�3��/跾6"s�֘&�"[6��ͷ$0�#A~zt}k#�����,��
,���FQ�o,�|��~�=��E �(HS�O�;xQ�;&� H��Rf����n$69�S�W�����,5�xA�}(�3�J���i��Y{���������@��TnIѣ�M߻������%�L��U��Cn�r�щلS#2 ��K�t?t��xb��Z�zn��*:�ߋj���%5��O�zv�?�L"D��s�1v�Br��|�V���<�[W;�$��fh6b�t
� ��n)ބ7���^^�SQ�$0�Ѥ�Xfc|IV�6�w�ךX�Sc|���-7��FQ�����$�?�OS8P������:�qސVчsr��יc�$��n�۟�x�����h�$p���%�Sm`�����p\�I�{��X��-K֐F>���L~�v��F:P�H��'�KG���S���j�|Cr��^��!<6ᖥ)�*��(�8b�2�K�˩﯇�l�W����Y�û��џ��r� �~4�HkpŏEql=�U!#_�t��DY "}O��G�QW�P׾�/��_d\$��n=b�������·�z��2�6xLv�q��c'�p��}h� �URW	� �L�g�}�r���h��k���i@�2��`�}���4߾!Cr�1�l^��&J�7��znz%-	�D.��|�P�@�������t�P�dv�����oV�GƱ�٨�|u"�n�j}b�Bu�}~#p�K��jm���ϣp�v��8��H-H���!OS�Wx�u��\s)���\� ���|	 o����	�^k��KF�@���6q�D-�$��eZ'P���ӽ�oN���wl�y�cTi!:=�̻����'�)T?�S��UZ���_=�i@m����C1�Ā[�o��j��zB87�y� o���8@� �N��f��/:��� p-#���ԕ�A=&r ���^��a�h��ى��>}\6`Ջ�3��T�ѧ#o���Lb��t�m��s��a��>��!"�����푂j��!$��8b���R4Go���Xd���>ˑlMȾH%y^-������PB��]�4�v�M>]�r;�[N��
��D
�_�/����8V�GIdR�_�����_i��z1�����Sj�)�d9m��g�uK	@����i����O԰8���/m��}pAfN]�D2���`�<3��0s�'����D�W�]O��=愯��P�y��B���=���9�
J��8'���_?\�d�lD�n�>�s�6X��V�(:~/йa��Fz<��E!gD�-l4"��K�^<"&��a6�Ń+֜�yC1`o�>�X�A��eR��� �����X.�DQ�'/�\!ї�lT�Ձ�t�����2�����3��,�!��n�7������z9�ІR.#2��M������T_�O������/T�>zҾ�ԛ��O1K鉳�/�K�:���epJ���}fQ�}r:����'��C��]S$�b�L�k�v	H310����x�j�k0�������Ŝ:�j� u�!��8g^��I���޸�#���=�L����]J���>ռ��A�}��'Y�x�}����2�j��vLV�f�>r�Y;�@	X��v�����*�;�7��pQ���8x����A����@�����z�m58�b�(&���/���#���)��R�bN��W���GΙLh�!�Y�dG����J>��Y�>(��Q`�lB7�o�@(�c�I2]E�����i���Ѫ��� y�j��ެokY���� #��g*�I�w���!����c��G���̏�;4o�U������ߖ7�%T��$2�)s.��iV �2�	�U�X�ڽ�s&%�ycw��
�٦�����)N����",`���Y� ���Ç0��O���`BbziX' �O-���s�r�z@^��I(�}�b�Y�{������Z��n;������������Q�@��u�jލ��S3��k$�|f7��O�N�ԬA6E**�@�L��y��[����H���r��v;�%44�u�����*J�9Ar�k��� 1��50��4D��:�5EC9�? yVd�������󰼏�攂����Y���q#?��t�yTzX��}��Q ���w��5(�(��פq1�>0�Cz�A�@m*z-�4Y���M۾�;!;Ae��w���+�a~
T�\�>}Pt�/g��m���xlE�õ'z}�/�������/辧���~�m��?WWW�ތ�m�w_SS�Z}
�� ��,�!e�h	[Y[[���q�'�NGӿ��+� ykop����K'�-��/B�g��Gį��?�4���[|g�K6Hk��+��R�vw/��IU��T��󪯍��7�,�?8h5��x~@X%;���:���E��f���E�ˁ��g�i�A.�������;6�m^�3��j!�պ�;0M��h��<�Ա$���|>������Z��am�y�i�:���<�m'���g�P�D���� Ô���olj�A0�H����)��q�c����Q\O�T��y��"�-�q�ыb�e�!�����+.��Mp�q�~Ȱq�D���� Iz.lؑ��u��O7����?��"!~�i�d|���PD��+7�=�C?ޛVN�2�y��sڋ5��:{�s\?�v���hF�?��ņ�� {�o�#;�RDy<�T[~^"�'���D�����m�'�d�_�0�-w,�_�
��t͡Ob���ԇ��%��mT�y'�T�vBxr9��o��x1�rD$���Q�|�^r������YxX5/q��L�mw��gd��{�[�)+���:�K����m�� �{g-h���#�jt��&y�G#�Fr8z�OH]��%���&��{&/��5"y�n!zU�
�4������l�e���kt�F�a(����^��]���X'�F�"������zg��ϑ���¶� ;0�i ���l��7������B�ut�xj��|��Z�ri~�Tw�q�ȴl�?����B����ﳱG:�<u�KWr��w6��L�eu�4� ��Ų����F^���-+01�J���
��%�o���(N��7M��U�&�v�D��˷�J!z2Y�d^L���O��5�ہII�!m
9���_,��&S�J9,�R����U��<��`���gb���D���r)�_[S����t��)�\��N�i�to�>�\	��+���@���L�uJ�r=C��2%�M���GB�}Z����ON	+E8���5^���|����N�*ec�ôLW<���xu?����s\����_B[t���K'{2���-N]�opSc�&Q�whk����bg>��O��V�o�.�K5��ߘo��Gq�$�Z�g;_T�@�;:^'�'��.O�B[�
Lr�pЅ7,W�f�K��w�.N�!!!���y|�i�:��0~��x�4'E�-��=�]�j���c�����?��,��%B=����#��&�7H��D�,��S|�Esu��<����]i:���#L�n�Â�c����֛�Ė�P���ٮ���L�>
L�M�ypAb�\�zO�����_��y���o�E�趎�`�R����;�M+�c����e`8�k�C�Y^���bb����fy_��Euê�f˭�fD�ڵ�`NN8-���̱^G6M���RH���<<�&�ߺ�9R+�p���x���r~RRRR+@�=o{��{��&#Q
|#�p�������A'��2�T�����L���"�dN/�>�Mk�-�K"��F�9��>}m*YjC��y�ɱ�)G���%V��ǚo|��Q��M�4���3��q�_��9+)��$7��QRJ������}�I����JGTX _^PJ������#k�Xy&�BJm�x��LJ�	m��,t�Ud��,�����ʘ�-$ե��ñp���g'/�:sh_���Dr��T��3�"._�HF]��y�.�����r~S)F����2dv�E��jǫ��xyӒ��R+3�h�:���B��Uz3�,����MŘ��ϓ�-��������%�����8B�h�e�G�(��GFFJZ���
�U��e�g��L��x���y��Gޑ�AW�˷K>��kQ���FN6�ˆ橉	��Poy�b��e�=�rg�*Js���J�6��U�7���ie8$29?lM��ȧ~�T����3�
Wn�%Rs���l�WbҔ��f��?ۓ�p?����5tJ�����et]��k�R��b�?�b0Sm `�K�n���������f]%��ײVb���� ���Ã~�8Jq��<R��ݤ��Dy���@ҕt�~���GQ�h���u��@}���k���::Tg -�'�RA�-�$���s��f�|I~�K�k�*�iz�S�{�j�������݃��BN�ܫ�AEh�?�z|��un��� ݣ�l�V��ǈ�I&9�<�և'1�gKn�.a_�����P�f8���;!�V�bűtBBB/hB��O�r;���%k٘������#Jma�� �e������B˜��&Lb�?o!��9��"_�3���a4Ddr�K��I���~�V�㮿_�i2��d��D�j��`�QD"����WUj-�a,��<��r��o�Q�k[�e�ӗHN"�Q4?ɸ�썃��Y�i�톈�F���������k��_�~w߭2ǭ�J\���V�'�7����3yj�I����0�*�ɬ������BA��,Qo�01cCfm]���4g'P{�a�+Lj�Ru&���.U�mԢM�:T��^�[`���?�;ȴ��:��A�b.�}�*=pn潜����>Y %J�Vy��/jr\�?i?C���:��20Ni���$-�Ǚ@T%�AEU��i����{�Q*���{4:%ؒ.����l��T���J�����)|��(������O2�y?0/�آ���n8o��*Af�	?R�h1>�K]��9�zE��A`�_���==I����
��F�h\s��F�Z�h᥆[,ʐ�����2d�8���1����M���@���I�"~oO^q<�P�x>���&���^�]U?R)x�Ƶ,l�Cj��� ��k�N3D_El��"j~�+Hq���1�mh��}@����V6�M*c�Uy�u����R��nȵ������{~]�+���5ȏէ���K�z0HT��$��Gq��.VV�Q���}<? �|�_C�/����@��^���I����v�X�<���UsL\.d�{��kC�l*���q,�+�rsM��Y�?�,)��V��iщ#i�Z�m:c�c�V����7��,�7�v��Y�)�3D۹��i}����	����H��Hk�9�}i�q��[}�ij��p6�"����m,�~��E�2t���Mq �8��<�'#�Q%�0:x=�����V�Q)6�I�u�g�l#r?|�`�g=�:uAS'w_��vH�KRp"�p�˰���=JxD`;`rɆ6|�%|,��fd�[�:�0mHDrE�v#��$Ve�l0������ڇ���r��pR:�I��1�2�Gb�7���uaaB+�Y�L�o\����91a5�{�%w�ӛ�鄙���ܠz�4'�;H�̑�T�	��\X�I�e)��8���2�w�,/��tk��A�<�B#�\�q����5�T�`�@w1��2�qJ�����`q�_[G�O~V�$0V�w�/Ps�h���[C��v�X�o(�Mj�HP�
��]ё�G�o\_�R1���i��0��Q�	���%��kf��9L\\5���a��K�e�!� ���m��s�ꛁ�'�Q��q1D��9,���F�{kz��
�>�2��F��a�
���%��009�� !�j��ݱ�a���q�\
�Qy+1=��2V����:�X���ku�-�hizf�n�m�#~� ����YEf���&^���
�J�˪����/9SD�M�'��������᜘�_g���J����j�ۇ����_Ә���N�\�K2قT�iE$M�����-���g5^�F}CՏ=�'ċ�A��ƨkW[�4[��HF-���B�|R1l��\�e�p��>���v���gY�iD���4qfRU�LP��}A���l�A}�`�����c����UL�NCZ��aKs̕0�s%�.�2�`0�[,����&��>��\Ú�M#_�m�Q=K�9]zrUY�����T��(�CX�=ڃ ���d�W�	�(##��p��z�I��N��:=�1��h �(E$����ɩ�V�O?��&f�U��"++R�`�jȯ⊂e���V�� �t�AL3�F6ra��0��"��ԧ��-~(>����99IY�z�
V/|��J�k̈́:��S���ܧ[����5��~͌=/�aPf�P�M�Mb--e��B�ߊ��5P�r]��e����N�l�hW��,�7�8$��r+���𦢸�������D�01\2戮4�)�|&�r_à+$�2v�E�_�#f.�x�F�E��o��P����^�1�d`���DGv�]ܽT�
�Ó	���ބ�1���@R6�j��^~}��CPP��m|E��$�֥Qe�:�)1����g�A�2	˾τ��E 7<��{~�K�W�-ş=���4�[�RPZ����1%�"RuFx>�$t����ۂ�aX,��?> �**�"��^��Ҡ�=��5�k�?�2���^jm9gT��[�ك�,\��e���ќ6�C�L���NH�g�;�G����A����|H
�6��_�2���1Bh���0�WXu�?�t��2��Qf/\�n�%�� U��Q�BJ��`Fm*� ˿���bP��w��S�Yݛ`&����Fu;��sjD�X����z\�:vu��|N0�1mucj��C�q�����u,�m	ም�^~v]޽sl�>�v�/���y�=J0�q+E�s�(�}w5�;��=�c�G����������(-ً�
�;mV���
��.�٩Gk� ����@I_��<�i�4	��uT���"�E�p�0��}R� ��u?�L.�|�L���n��J�%�yD��	g�����W���%�m)��$M�ʓ�n;��?ئ)q�5��+���P�Y�kb���J�,���׼�&�{�m����;~cKnx�J~��-�*���#��\��>�:�f0M֫Y(Y�;ϲ9����d����#lu��kO�+��r~i�^��0� Q�V2y��4ۓ��ia����T��yok}ߦ%l����"�n�g��n��k:~�dQ6�u�Ifa�3��)9�! �l��Ԋw��f%����cэ�pgp���}����֊i���iCkRb�@�uN�w�"J�-���hi�����z�+�֢�5\v��IE�ņO9[�\��g��Ζq����r!����$ɠ�|��';��������������B��K�܊�6!�Җ�IJ�/W4'/��� '2Q�\e�ַNN�!������U�'����i�Qͻz�Ŧ������v����4\�a]��ק̘^aN�Ou�����ڨ=ja�?��}�������+N7/����XD[4$Ǫ�}�c�Ȋt>�1�o̖L�g�m���Ee��I��Di/�`�jx�S��4�B7b?�C���h$�E��6� ��N��@�-:�ӀH1��:���f
�7+j��Q�h�Y��TwR��5��L��99�����?i �&)/��arE�נ�X�ts�4H�a�U�&b�N�~�5O�`5�\��(�_&׬\,נ\���� d�Y���Q�����9�O�H����_�z6����o�ˤG��9:C[�'W��dV#=��ӯ�D ���.���(~% �ly��]/I-�z�K�����$��rs�i5Zȅ
>�._�N�<��驕��sz#Q`�eť�[;x0;k?�XU6�F�X4��=�\��X��To��.F��뱊�:�a���s��$T���3
��ZG�2`�sXW33�bf�5E"�Rk�?�˕;C�^2�j*��{g�����\��rr>$x��� ���8J5:�/����17�gW1@���5�Cz]��x�y�l_��ޅ��e�hw�?��bA�7�{�,�
 i:[B��x+������@��>��xl�N��;k�d���]i���,<����3��������Oެ�;��x�T�F���)���x	N[�eQ�{�w������Hr��\|�Ԛɿ��1j��F���f��k��[.'ʽ��1;PP�nRj	&}��S	I�!�cIk����t�+;*P�`,�}=��(�u��A�Nz�촫ꋮ���c�'d�NrW�\w�{;��U9v\�+�$6	�N���Ym���	�B<7�(�}�aj#2�2��4���e5C�\����"������)ݚF� C��~i"z)��q��]�����F3�t�� �SV g!,t����Z�[�Aտ�ӽ�����c?@Z,�I�����,�B��Y��,o�'"�u�l��;��n�?č�ٜ������'NH�X�eՙ�׼L;�e��v4j����1
.�AޗbB8�3�||���C<gA9U���;��2ۭ�'����y��N�=�p�Ev��os9�{U�8��m��	��Gz��=z��^��1I�!�ar渚�.�߂bI�9ڋ;!6�*k���Bu6���n�`�M�$#�i5v���}a���������:%��e��?ܭ">h�!����S��H0�#-��LL	��h�������l�}���5��ef�vC�0Et7�C}|��{� Λ��J���4��[�@�y�ˠ���"��#���TT���r��=�������x(��Mʞ�H!�0!$c��lI��d��c�����al��oٷ�uEBCv�dK����}����'3c<����9�u�u�	�4�z�#K�V;�Ahեn�t��w��+Y~~���b��������Snc#�����/B�ܿ;�Gu~�D�PVXtJh�]�Ƙ���v���ތԴ/:&F��$�U���I�ŹEEf$*�Ȉ��b�RE�X�0�7+Ы[��� hݱ�,�'�_h��4�I���tfv�����$;���67ֈe�~nKz\A��m�gq�V����V\���?��)z��g��\-�?f����p�G�_~8u;ф�E#�.
�j5j���{��g��gYߓY��t���5�!��� ��{s����p����$�+F�l�)K�N�̳	,	s�_j��v^���/���� J�Ϫ׺/�U4�"��$t>h(�����.��6j����m��d��� K�� �2��̚��|��I)3e�􅩝��+q�o�|�-d��x3Vh�=voubS�;R$دnOK��2�LQ]S�5A��ϒɯ<�8翙>�(#*�#
���]��k�S��9�BI:�VW_�n�뽠����㴻�TL��t=��.	�'0^ý�ɫ�0��-cǴ��ƭ��=)�x��s٠��h��7B���n>^#�&�n�?U���GI-Tv!  �jJ��wǔ`6A��T�{��k�rq4'�����4�]��[1��{�M�J;�;5������D//Y�"fS<9a��Iܪ�<k�&_���y`�{/$!�=�T<ax�x<�:��v���zW_R��̣m�/ �X����%�'�`��I^�-�G�+.(��v��k�)ذY���ʰa��ǚ�3k*e���J1[4a��BA���l�2���}�g^�x|��k�D��PFd�UhXm���*�dO�ش����7C�"*�	�.GP+����k؏�Rg�y�,j�{�^�����g�P�B�nT�8��kۤNhOQv��ء�@v�N$��=�B�g!`T2�^����9���~ں��I����ډi��F0�̊����=;�S�w�^PB���7�ӯ]G%�&k޾�m��4E��IX�����/.r$�[(�����D5oBp�k�,Cۈ�f7�G�1s�����EɨHA��������!�w�Q���E���0C���jX������	����z<�	g��rA����B1��3,��m7i�`�X����-�̖����O��/{yr�-"3��z2��r~Ө�}3�B擿�>#E����d=����������"Q1���y�|{J*�D���рW�ֺ;.A���hT�nZQ��<깄��� ��K]��mEi��lP�\99��u��`�o�v����Lo��O��Y��K¨� �c*���z���T��:��d�+�e�,�py��h�%�{:���۟���B�3�d��g�����s�vWPm^t�2��n����J������T`�;&|�^��m�^q��f>3aB!���ԛ��-N)6Ƣ

��˔�>��Me%��~>CVè#�Q�̦P����e%��0�<.�jȻ��w=���m�h@ͦ�f%��{^9�IW��;gg��D�t�z%��B���w
w��f�%"�7�Qϋ�r���,������-�^5�_5'%��R��P�'x
�D����/ڠb�֌*�y����[[�w_�%�{��9�
&'�r�i'ѱ'�i����]{��%���(���;˨�L'��˦5Ų�I�q�6m�I�ѹ�����>=~��5Vs����oA�M�P>A�(���|��3k���1�WJt�Ӆ���l��jtP|���ZTt'Ug�`�8-K:f᾽=�%�;�z��f��N����W⋢�������t�V���W���G5�ʼ�O��5�H��rTZ�=���AU����s�x�l����$�80P��Ԟ�)EM]y�eqC�nunQ
J��ys�J0��y��x`���e8�~9���Q����hxLuRE�%�]��+�������X�,��E������fz⸝R[�e`����|�'?&�ӳ��6���,>���
/<�p�A������K��ʏ��D�$F�������������yէ�`��mO��g�d��os-5� N��4���/+����"�6<��fk�Ʋ��Ǽh���e^�8�y�i`{�RO�����hP�{��U��Vv�:nA����<�B��^(+x��Lг��!�G���W�.ېs���7�բo>~�8�������O�BP��0��;�
4eOVᄷ�j�-��p�Ohɤ���/M
Ui��ŒݓS<2����{�mg��T�-m?Æ��UC��8kl@��7V0���v7�k���ג����Zs�8��Zw�&7Mf��57|��LY�k��捤��=A��1���L�:!I�󨉂��5�JMgkgGv�2l�a/���[��~w�0f���W�` jq�5b���A��\�&�)vy���f�([z#����)S��lV	T��sMƯ�NY���k/ �ah�n.n����}�	%pV��h��&N�]���+4�l�Ɇ`�y	��Z�&��)�O'#�������	�V�y����+��t���3&�����v���p�������>Ē.ߛ~�Y,a��?�ĒU۹2aߎ��蕛�&(X�Z�L��IU��>�/�e���H��e`Zz��\_Y��	 �;�(���@u�ߧ_����k[3v)�ZW�_e�!��鸍|8=����S�Ƈ��2C�V�>h!��S��u�����ü{=8��Q+գ�/�}�PA>�ꣵEV�Z������%#�IG�=u�������dU�'��d��;�7� o�P7��65�љN^�:)�w�B�ŋr
��**\Eї���K����yH�4z07ː��=�{��2S{��<O֠�����W��rq☩��IsR��U����p (�=$lﰽ���$K�;��ו6˧j��T�UX
^sz@�I���b�q��#�S�=�^���mgk�����\�!/��ۿC8R����	��/1B�ZYY��7`��\��S5IXDboh�� {��鶞r��[K�տ�`W��k�Q�<��4{Gڎg�:[�����]}jFZ��e��W}��A]�J��PM�9���${���`��	��hWl�Y��u�w��e�b��'5+싡'kߛ����[V�?ι�z�
��s}D��Ӧx�h�,Nj=]��VI�bb<9C��m������!�n�/n�R�;T�^yj�>#
���z�#^��Y���D��F�H?�j���9���1%
͆`�#:�:$]\��Z�d��;�1tJ o+f�ٸ�a���P��|G��r��c� ��������g�3��酔{��K`a/0�f�N�Fff�0�[_*�Θ�eD���\T[��I�Z�����nX7G�*8��Yb`���Ғ�2L���a�8 ������Ҥ�r"؃C�hKY�K�D0l�]����3��*L.��7Y�9|����~D_���7�]�g�%�$δ7��62�Cr��Z[��M{5�Om�4��Kǯ��eM�2�%�Zp�^��� ��Ï�<��[�4ɱ���-���i�	O �|���i��6�ɫ�Ey��Ѣ�����VN`*�+��5����5^e�u�Ǥ����R�Kw��?�)Ľ�g�|�4��f�\9:�\q��NI�z��	*J�3~kGP8�,��V�8J^C{�G8TE^K�B����z������m��He���I}�{x��P�a�JQ�n�D���ԑ7�h�%��d�8�t?���z�S��[�mo�����9��{x�BXy�2�z6���*
�JHHxԂ7ZW��d `�c��:�W��g�>��i��C��	�<��Y�$��)�8�b	��Pa�MD��-+y.����i$�JL��#���4mBeMC�H��'5��G�$����Ɯ��?S�������[cJ2ȈP%N��x��Hׇ�8�a	CR|�%l�:�:r����]ra���FaW���^{��@�:�%��#?������j�s	��,ȞC�s�aF�|$�1���&����_���N��Υ3�mmm�)�_������JTR��=v��LAǔ%��C��ݓ�k+� Q/H�:���G�n��ܕ�N^:�P����ܬp6x<��)��ӧOi�����R���-�H�	�C��I� ��*Q���PF��x��P�,�g>���*�I�n�A�Ւ �~TQ��������˒�Q��W�n�kF���c�\c�y\�^��Y���N���6��g������/�;�$K�A�p��E#�7�x����4��W/i���r�^Fy.n̲9]RU�+�c������S�")I
+�RIDZ�~}oơ��s/�,��V��$��� �-nF<�<7�*�&�/ٍ�}y̯�/6��@�Z#�BU���l�lb`�K�(]���E+_����w^��lL/�����g�5�����
�.O�MS�y��]�Z��ͯ5\�����!��b\e.u�#ЎpWXC��@��J��i�� ��?�5�01-��K=\A{1ܰuo$3D��?p��=Fw�؈%�E���s_&Դ�k��k9x�%��(�x�[� ؐ��Z�5/,bu�Ă�x��M�Њ5���O���Tg������}~����@�=���Wj$+�m���ޢ?9���)�4�%�*kX���{H����'s�Q����v�E867���<}ݟ!�ۋ��қ�'d��GJJM,5�GV���BSt���;gOD�&!�y��R�0"��P�1���i�n�*,��;��/�c~B��L�N���{�%	��Wt�A�e�i�ԑ��ډ��i�����̿�\�u�'?���C�$�tqFZ<�vXt����s�p]��8����B�ߊ�]�������`@CM0IWp�Ǹ���G��=3
�E��'6��l��.i��탗�l AO�s�1��X&^qHN�w�;rsKJ&&�o-�����#D��߿ed�[W*t`:�v?L&�5�/�٧��:��7��l����,D����U�%"��V�/c�SSS��F�[���N�5��W}`�~�2Gi�c��p���LA�,��<�3^�<ۇCů��aS�sS��K\-䅡����9/:�s�b�EC�|40�||�Zj��]a��]|��{�P���x���s_u�Ƈ���(F���/��+Ӆ�x��4w����E�����S���+���
�Jj��!��:�[���?�}��ՏŶw�� ��M\uѝFqIX��̠8B$���-��ƍ-=H�$�+��O.�N�`fCeT��`�x�ƶ�ԯ�P��J��1�'؀�J�I�g�"L,���99�9�n�4�ح����!���Z=�d1���;����$�7���U�)�|.N�.]���O��u�me�m�88�W9����c�U�x>m'ժgO����O~6�a�%��p����ӪJ���<�#$�ϥ$�����&=���w�=͍LLd�m�q���G����N�zE�}��J�f�h�
'�[����&%�N�vo�Duީ�����o�ߨq59f��� �'����H��<�gS��*���#^�ߛ|�Y�="��J��CJ*��r����N���,{TghKG��C$�`g��c�1����Pe�{������������r��D � _{<��*Y��7��Xy���M���-�SaJ�`�pC'3~��
`Wϋ�-1MF�;2	&�c�Q�,q���q� 0���HWַ�oV~X�/4^X��~��. �[�J��̈́oH�o�@����,p�d~�6�xw,�#������P�!����>c1�_�"G<���~��ob���HC ��wk�\L6wk���JJ,{������(�W}��~XGxĜ�,�<ʌok�D�q�#�u=k�Jo�#le(LV���F~m��N;We���R,�bµ-&���>�X�I�W��b���>�;�H�t�Uћ/օ��P�8� �m��&�m�����\qA�z�]F�{n4h ��O�Ozjbз�Q� �Z��y�Փ��"'��و�j��Ӵ� ��r�e�7��&b �p�t�+���i�����M���:E����s)��ΥWQ�N�������˞����
̙<�沺��`�a�]���:.�XD��vǢ���Ew���{��l�p���d?�{�K;���=́!g�T�M�/�/��{d�+Gg
�hyX}�<���;���<��~~M|�E#�H�xX	'��������6��Z�s/��JCW����BFx�v�ăl��Ċ�>�����#߯*��A�H���Y;���s����݃h}5�VT�A�K�p�ܦ�w�a����&�����h���鍁�ӻ��2��G�UP"�6���٭�q�s>�bh4\9��v�J9Ӧ��_ˑѰ����G>�*���.dz#�zn5@�J2aLkm�0[p���5��[S�@�����z-�8�2��.���]5����7Oqw�懓$3z���z�3Ur���Z ͦ�����;D��t��ܾ};*[��xXF�Y՗�����a2��>�5��"{�4�gʲ*+�H��;���_k��?\�-~y�A6-q���|���y���.8k%w��'B�#�2S�`�j���ŭ�hT=�7Q�7������eUOX�6��7�~\k�_�N�4�N���XS�^��l�����s�� �Cv�(�4��K�]VB��a�?��ʟ��<}���p���l��i�뛋��
�]bK�3�Wc�>|�:t��\^~������m�p�v���4�R���}^�)��)5:Le���,Q�J�3��=�f�� ��0���p׃�,�վ���nS�MU������&��TN��0i�嶂��m���ֈ�-���/�b��qOn`�N$���>���w����޼�$��]cϯ_��
������ju���3�bb��O_딶���bT~I 	�=#��|U�]V����g�|4K����ܺ�R����Ur5�*���ܜV�eAS�
��5&&�}l���Ob�4D�>$��偡�c��N @������<��V��z����];O����'}!GgV�fͣ4�%A;�%aAK�d���ᗽ֡E�s߅�"��&gB�NZջ�NtB/5--����3��(�Y���Ͻx�N�q���&|ML�ě7o��mvL
�[kN):E��0��>*qZs�W;�����dm�̈7�r9�����Sm/Pn/$�ٓwW~�9��u�����(��v��-$�?0i�l���䯉����owz��
�PR��_���'n�i�jr�rZn�&X�	 �L���PਐoBOe�m�����>���j���^��Jf,	ra!�݂3Df�N+}5�~_#����X�������}h՛7e�� \,1�m�i��	��8mr���<E�����ݾ21�l/����������Q�9��k]�'xG�����J�Qϙ/w�*�������B$���i��.��H�w\��H'U��u ȫ��y��_0��Gk�%�@5��̛���B�ɽ+���<Lտ����w*X��&���ϗ~M62ǰ"����ѡ
��o�1�p�;�v<�Zq�AƐ��5�ܷ���7�N�d>�$����%��&M֩�j�|����Sm�9���jlEg�h N*�u!����xdAҺ�)�4JCC�F��kg٪MN;T��/0i�{��+-_�d�.@�/��s)׬��?�ֱ�!����&��W�1sA6�A'�26���u�c�����%�G:b�to��Z�R(a-�Y��-��	(�`�
yKK��������ۍ�"�����J�&g�^�x���;D9�1��q�7�UY��'G%����G��J�e>�)�8zC������f�Piʰ�ZZ%��ԑ��&��[J�՜n(��K���8��b�Hy�1��<�5!"X�c�P*�rX#A�v�Uf&i����[߭�E�ߍ8<"�q8�G~x��'_+�����:��Q���9�ɲ#�t6pm%$�0�e#��@,K�G��Go*�(�h"�r��t�Q%�2���z]&ɼ��8�Ckwg>�,�X=�m��;G��S��¯���g}cՔ�S@C+�0�i a�;�"�}���5�(�էh��Ѝ7)�t�������``f�3s������ޫSO��S��1b��X��n�պ\�l��9������L.�!�)��-�a8��6ZP����N��i"n�x��e�?�7��rI����H���h�zމ�W~����ow ��1�b|vr3�%�^���+k��W+���&5���]�������Kx#w`Lzu̴UV%�7)�C�/�-��e���Q���lwJ5���߿�I��a����C9�^��f��t��M��K��.���K��ƿ�������gatU+�Z�k�)�K�L3��Q�J#�\�C��@a}�)����V�ky.����m�����V̄k������A�����黺�L�:T��.�� ���օ�|�Y^���Ц��Id<��祜O&�0e.D-h�yV��La1�#��qj	]1�y*fԕ3�0^�[N�f�N��w��<e��V�yۻϗe�ֽ������ ���˰	�ē��/������z��� ў/Ǘ����m����L�
R@U�T����D"���h���)7D��ᩫT����r��q�΄5��́����
�_��MUR��z�f�{�?C`���Ps�������}�}C:�*�QU�w��w��#6��*�9��g�-8%�2P�8���LS���D���p[ܥ��	7�����14� <P�/�)������i�t0�4!�}��*YLµ���!)�nR��vŜY94Z�P����>�7�?9�	�S�C�jF]��4:���bGU��?��3�s'n���^�vT��h���8EM��%}�M1�� ���V�V!kV��o�py5%���Ѽ��jy���"B'�	'z�ʌo��V�`���PBv�gi�W�E��.�u,}���M��ʇi_�~hikSj]R}��J�[��*lJ��\Mq�#ߒ���I����
�yV���'�g�P��%�����*1�WQ�bHG��?��eb�O��(~q�/,.��k����%l��Ύ��M�}�z��#:����͡&��˭��Dtdz�eX1611���~[���������T�ݷ��x&:����Ϯ6)�#������M���-C��qg���Z
AV�!���+���i0���F�s��}UC���
I�R'�g*�j�:M�w�k��������Q���,����6e��먹w[[Y}m���dzXgg�����k:'��r�������ẗ́�'+e>�^k1T����A}+�O��0*�E&����ܻkT�l�v|F%�|�������H��UX��&��i�@��jO���X��E��LήC��8̣��8��ז�*����i	cj��Ԩ�|��7��cZW��Q�|'�e��������cQ7��T=����p9�������Y�+JR�pUT�m�[�ɷ�±����(l����;���yE���G�a�g�W	��(�J
*���6��7v��R�Z�Ǩ{"�� �j�67�c�:����żS��#���}���9�!*]��/w��:��:C\��"�ޤ�T���3=�}�4����ѯ���5$DP'�{�N�T�u�8Ai�TL�b= ����
sR4�����M��ϡ'?���|��?j>�k�0����nNpS�����DH�bٞ@����Űɘ�'����2�x���k�\���o|���V�x���H��F�>>>~��mx�TTT�Q�lFUE�a��� ����p�Qr�Wk&L�Se��#���&��k�Ȓ��`p���
��|�wc��G���T��p�>�O��,�a�P����;��\BB!�$�"N7���5�z%���b�gP��=�n�Ĳ#2"�Q�0�3����o���˛�6`����c��}Ht�Ć<X`�E���0$v���Gd�sIK6�����j����!<�������Ω���JD��F��^X9�E}��x̉$w�7�������w�Ps�FP��x�-G2����3pQ�^t?S32���ʱ�R=�Y�ׅ�����Q��"��S茐�)$[r%��談�ڧe�����{�Gzp���i�IO�ҏ�\r�����8�_z�Y����3�× ��3@�-�R. h����)#"hhj��pcg�zR olV�1��-r�Ӱu�q���B�1�v��[#D;���כ9tE�r���l,ʌjf~�V3+���A�=��yT4��ѡ���~�gΎ6뉪�G
2��4�[���_���Y�G��b`z��l�i(�=\��?��j���s���u���h\�UB��8�Q5��
�>�}��Q 
�g���1UaE�=�W�hN!&�$���T�<oG���Q��iu���I�2�>4��,Zt�'镳P?�X�h�h���Ee�hr"�_Ư�����]�閙�Ow�5��q0���b��K�z��x]��2��H�-n��#@uK�]d��b5 �6X��Xtkdv���N��� ��k���L��E��¢��Ƶ�t�ij���v�%����h�ԗö́�j·��������䁢�7����� oW ^��w�@����2]���%"#�;x$G��9ұ���J���,�@����:�ô�����U���|�Zd��c2L%bQ��E���h�:�Yꙉ��E�>�3f�+S���e�z3�a���#^���2=�-e���%dz~����Ml��sl1S\�x�x*΍��G9�Z�0{��t
�\�tp�_������������ ��هN�{�4l,Ȉ�a�E��������X`��[�nܸ�A��S$���z|&�i��8K��"�T�$�)��0O��	����Jsވ���(����:ޙ[OY��o����J���;�����b�|���'�,z.�񜩚�==jÒ��bɆؑ2�O,,!<]��3r��eM3I�N8�7���&V]k��r�%��Pp8�&����p��g�&f�g5X[*�Q�%��*�ee ����M��)ӣ~f�k��J\q�&��J9DvX�0{�09ejf��8?��x4�f���Oț�r���/8"��)��=�_M�$�;�F��f�o�R�G�Llן���D����±���Աܨ4##�N��}<6C+���L	il��='*)�7�z2@DO��n�%8�[�+��BO�H%k������ Q�g��2,�<�$i7,!`G�[������V줪��eL_O#F������5����:/��}��oy���3I�� ����ݛ�`��n��+ԧO��\�a�T��}�^���3���󸚰��۶Ww���'=Ha�73��j����%NOe�`ܯ�z�caٰ\&e4U�|�	�h
�����\t��`�;u��n��|9`+���gT�.m��&!q���[(a��v�|��%xMZ����3J9t�\q�$tߪ߼LZ��ÜlX�͍u�%��dl�\C��ݙRV����b�-����#_1�����b.���,�YU�i���7�o�����>�o_z���H�А�V���_z�����#%��=⃲[{��@�	�'/���j_���If{kpJ�|���X����!�4���f؟��u�������t�a���/���n���;����9��H��T�6�6I�:D?xN^%�<��CO��5�>ZW��,x�j�@OPG0��T�Qq����l�$�a�t6"�./�N�uT�d��F��=80 h)�v8�ȏ�,E�5�j۰��0>�"�+�!�;2(��:��6^Ev��z��H<�hf�e ���>I)_w�Z������V厧n����U�k�X��b�\W�.��I��z�_N*����A�yAD���I�h�AQ	��4!�w�4yZ~ۅ����22�:"h��쌙�;� �d�ib#J����bȻ��A*��޽���c�.��	K~� ?v	y�iM��
!a8H���H�bB�C���;���}pd'�u錿��vQ�He.xh1ɗ�#m:��1+k~4*��v|�b�����B���]�A������ݻw�ZkMk��d�o?�b�:����g�������g��N��l�9Y�ѣ�X��b���5��Y4\�J~lFJ��
G!�Q�+� �!�m�����dQ4B��Z�¹
�,oE�+V�o�>Pea�"*//��,���s�|�ġ��X� �<�P���t8'e�~u�0#�R�&q�Ԩg^n��q��W�����O����10 t���9wdVb���smJo�g1c}=<�/���{�#�`�z�@`��7���E��Έ��ݺ�u�'��5�}[;;ã��]�x���yPl ���A7Y0G�$�2Ip���}���x�_��~}5G���}����-�Ͼ�"���íQT�a��c��ֽ�w9r��.]����I��;�RM������p���pb�O,������IR��].����7f@�<��ې�VE&�(!������E,�DG�i� ������/���S�Jw����H6�����x� >L(�n�]�8~N�XZ�/�^eG��7�iB�c��¬� ����|{3o?V�j�z�@b"�Iae5y����5GY��hFE��ϔ��n����-o�'�w�;e��˼ɠ�9�]��.i����zw�����<F��N�/��@4�@+[�v�/�]�@�"�:VL�)Ho�d��y	m��:��ѥ��O��)�`�,ƈ�/������]y���T��6T�vL��-p��:Y��=�d���l�]��d(��_!>�k��^�E�;3p}�/����G�,�GHCSަL�#�WZ���L��������b-�����00]��7�i^��''�a}(�n��˦�Q��xmBD�K�!��+��XMj�K�Y��A;d\,���Mq$�,��v��V����պ�~9�X�rẻ�g6�/�Y�:�r��t�W�Oj�#��)���|�ɵ����a�3���y�1��hbd�Z@�u^��k�O�,p��g��b� Ogo�X��~�%l3�Z"�DR����Ԥdq|j�f%��S'�n��{1����t,s�ö�<&�kx9�ݢk�+.�8A,쇓��y�0���ς�c��<X��g\1���ɩ�xa�V�_�����e������?�V��;[e�O4맃���*
D��`S��(��kUa4�*��k?2 ���~���4�5��=>M��m܀�vX��0��{��XB둠D߂�0EL�j���	w�����'�~�V�1�����p��Ta��A;ט���M1�9��T�T�]�����K����|1x��z(mv(r~��+@��ƪ�y�ECr����[4Ԝ��M�x�|պ݅���mpPe;�9:A��,�x�8r����/q��~n�-'���ٯ�Py�d�ng8�Ql��r��c�_�� �*�Z��ޏX�;C�tN*�J��)ꎇ~T���-���ۧ� �u-I�,|�������z�¼Uܰ%�9'�NOP]�
j^=O��ѥR�qM]�a}-m�/�b�&�d�<X�[L�IZU���ݯ�)s�[�W��.n�(y�jXv{o'y��>A��g"~�ڗ�fq���Ȣk�)fѲ���W���˴���U��?]i�	k=NȠ��}ڠ?���vS��c5��Q��Q�'4�wr}|p��&Źs/`�h��Ѝ>T���CQ9�f��z���ɝ<'�{�u�~G��e��$)�CA�����~�>'���I���BT��8���u��O$y�:`3&��ն�*�R5������m_8�
Nƴ|�0�ϼ]���<Zʭ�~Ik�#Nm��-tge��7�#��t���Ѓ#���ԭO2]�s��S<r5���}���j�Ϩ�B��i*�.�3-�dmڟ��07s�x�^=�H�qf����Vѽ�3�#��o��+��x���gRҾ�^.B�T�@��"����5U�/�4qSL�]�����qZ`��� �ܓ�-&WW��Z�vv��RE��4�+.�l��t@��o�O����ũ��"��2�������S�׳�*������_��>�'ܣ�����Dh�����I$b��x�ҭ�t)4�E�t�$\�7@]�%F �3�q�|�d�ݨ�s��8I��ε��lNhE�m��KnW�8(�;kh6#P�vo��},YnP"����T|����<LI����3}�R��r�A�V��۽�O���x�}��	U:��t�^O���]i8��!��O0,��W�����5����T�}K�ƺ:��ׁ�O1baa],�N�f�y�4��!���VG�W���0��ى�
�%������F�s��w̫��/�`�쳘�� �I#\��d''����f�!]�S
'd��V�m�z��fU�|�qS4pC(i6<h�ﾙ	�I��x2l�	]z��WQ,����V:�҃O�Ǘ#4Ի�X�`
e�~Ex���!T*�Lf/��������˱H]���c�;�+%ړ�� ��/?�MvZԼ�����SH��.�����l�m7��ց%7�ᒚ�XUU���������D�v7�>��В�h�-&xe��A~L�!]	"�9F��ͼ�V���g�#���f*�b� �o���%`3}�����
d����~8��`A�XOlT�M���j/���G;��Q/�I�.[�q�=�0=6z���y��A?�e|~O�����~ܸ�sn|�H��u,_�Y��������F׋�_��O���}O-��hqI�|�B�T�'ۼ��Z�R[��ݳj�7���*GEE����f.sr�ۓ��cb���#������uy���%��YZ�c=�`9��N)(:k�"�
F����E��\vg���+@[�\΢
�؎_Q��kԆ�����y�&��=oa8,�3��'�6��ɏ�h��NuX�gՔ��~��15L�Y@a5WB��4�����c'\�{}�{U�����R���z���T"��f�3G~��JM}
x%�p󟡫JzC����UPw��=�� AiUb�?��Zfh�0uA�oQ��5~�I��D�BK��5����I2$~f���e7��'p6�Ha�2�ߛXf8�7�H�#&���č�b�����E���'��(�g���G
J4�>K��+x-���w���`�!���	�Չ�f�<ݧв\5��]\2�A]���e��s��HkG_��6�Z+���!�����j�2b�0mu��+V�W��"ɨ;���]�?��H���z��L�z<Vs�_#٬��<8�z3��e�Z3�BT��#ܓ�����i8y%H��#����b�~�w����N�����?h�)������r�|�CLi=�e��y�g>�9cغw(ϣ�������WjF�	bɆ�2�"q������=d	�+U���j?�{�5�2�*dj2�ս��5i�o����7�m�i�&iF��mB/�>������
�������^@�M�#
�/)��� OH��-��W�x�F���-�/'VN �eO�eRBZ���y�|M�c݂3��
Oa��Ҳ�֗��N�5�-��Oq��J�~5��pk�F��G�������3Iq��h��su"0��+���z��Td�:����%��t.��q��r��w�џW�*��om��T �M/�\po�&��߫�»JQZ� ��T��6wsgw0������v��ݫ�4�ǣW�����^{�_]�	�������z�*�����.��W��]�<L7��i��Y�?T`����4bl�Ou`HJ�Ĩ���M+N.!��T�-���+w���ј��(�����|�U1B�کa	N�(�z3�����[J$)�1H�×�T����c(F=s̄C��2k��ǔ��{�4�Ov��
�e��3Lchpآ_�8%[t �,m��L���DVU�#m�R�� �{%D�D�fQN8��tD�u�;��BU��uh�N�|�l�Xe3��~I�D9���ȭd{�����<wg�	�TT���xT�/-���WGOA���/;F�U���q�W��gΑ~�ss�>�p����>e���ľ��A`*�������*^�K�\�9��(�B��-�����r�+=ܲ�}�>C,/��]�����?��e?}I���3Ń��.��=���A,�7Y/��>^W��ARvS~
�����i�C~�rsq@����Ħ�ĀɦM0G�w�Q6����=6��̩��+WZ�����t1�M��<�C�ŷo&�g#/=',8@�.;��ۇ*qB�{xxx7�X�Nv��b9�q�5�2�ӡ��+�w0b޷�5j��\�����}���u�eH�TE$�Y&
b�;��8����+3,#<�ݵ��:���{���E�ɀo�E܊�<4��hćc�R���f;�q�ami銬0�Hp>��=��������֤�I�l��Ř4LrNIIɏ���K�u�2����Ca<�Tߴe��j�zύ��d��Y1V�j�z���O��P4�6}	�ܸ�q�����]-=�Z��Jp!ټ��MQ����G�_"��^ Wu/����Ez�V�i��O�Qf������M���C������6����OR�R��+㱦�P\q��&}�-a��*`�6����e�u�[O\����$_����G��F^p�#�:>��#�%f=�x���SdVYII^�1;{���V�a��ǫ�k�2�t��1]��xt�.{�Ut/������A3a�2c0�|�*8���^��I�|��+?���E$Y�^LZ�y`���Zߥؤ6:dF�j����	����7;w�"^�"k]<"���L���z����ej��1)�U�N����4�F$�222~�û�,5%N�Tj�{;�z������R2�4�{-�����kW�&�Wvڙ[D��#'h�}��d�ۃs�V�T��~g�M�y~�Ut|��y1��7��9�C��a�dE�}1jvR&�S�,�ۮk�+��ǰgF__"�"ǭ!4?{lǒǐV��B_R��s��n���z7�M���#�G3.�PKR��ӹ��d���'��G��KG��J�K����t�
=��	��DGq�X)f�k�2�]k�7nX~K�M9�/)q��5}J
�[�)��#zh�^�p�Bp�r~^�1��Z�]k8I��J�m7�
~�o�y�'IU�����=Z�,����̕���]p�p.�������rrr�Ln3aöG��-��z�?�]\�-�hn�1�uw�8� �p\>~��6�p��~�X[|�\�ы�|���
����7w�>%6�z6T�l.U��N��v�24��S-O0���ẅ��6�繥de�fɱ�CZ�N�����'�N<x��t���y�J���^�Ԍ��(/�J��XM,�3p���~m=��/>�F�3�e�I]8<>+�c������ۈ��T:
b;�1����$Z;�Iehk�}��tE˱��u\ؗǲ�����������|R��ڍ6ڀO_6��uΜ���D}�7���q����v<�5�q�����LQE���ж~@��Rގ���s�(�3����g���)�o4�7`,Z[��8�H���o�;�\���h��-K[<^����z]P@T��L�w<���?.�%{����J��SfH�8d�MF��ބ���#;���$�de';|O���w��n�p����u�߯�u]�E�Tm���h�Hz�H��E�6oJAk��T�]}�۷e�d>�2'_�/SE
L��FUWW�����sd�	��b'~eK��N��#�8��% 3y�"��R1�*L�~g����nh��LM����TKPE�cei�r�c�𛼶���B8�L����D\�1���������[�v��q��%C]ݿ��?�i&�TNEA��wޑ{�=e������ ��R�!����0X��wۖp鎝���'�YC���w�l�^P'G���w�L�Ȍ��~��Ҩq?�vv����5�)�K���aY��x����� ��ne��1�5�r�,k$��s2v)V������{�������A�е�f��!}��e��gG�~}X'�b.�0���
�Eg���1ɓ�F<�ž<���	��u��(��?C��N���`��z��r�@�T�-b����~we?��_�Y��=�vB�u�5.I�0��"���UJ�p�zu����B��pW;2vz���	(t���~���=H1������w,,,�qɓ��"�5��Ȉ�1�Y 4����*����:�Y�������z�az�<�g˜$���t���C���P���¸|n�6�q�-5ъ��~��Z��<G/s��6JH�TaVn
�QU�( ���$��X��H�l�w��U���n��2���Q�Utt�4+>��A��Ŧ�s�d��а0A99�����3\�bҗ-�03w��YV�]ݹ¯� T�����7�^�=ުn��z�҈����z�	�.t�-�#��u��'�/��`ӳ%�i���5p���A�p��R\�r�V���}�E�8T�T�MV�!l�w��^�&e��4��߿G&&B�����Z?��	n�i�g�<���x��#�������T��N�j�����K����v��qaʪ_n�^z���Ty��5�S�)z��<$�������'�|!C��P�@3�q羬r@��\�Y�C,�;��ﶈ�̇n��J���G�"��ڏ���M`6X�����3Q��*&"2���ˋr�u���+Z=̦���?�짟���E��"��H*QQѷ�i8�$h�˱Yۻ�:<��g����F�2�����<�bD�=��TT��+�I=�doܜ���֖o��F�FM˷�t�ɱ1��F���݉��*2\�``��q�bn?[��ùPϵ�?�k�e�4�S2�b_�911�0�ӕ�1g�\�'2��Ge3U��B�V{�Z`l]��7b�U�xU�d���1W&�{�:�Jl�Uu2���J�ﳢtx�>PI��Ie�Df�ka�O�㪫��Oֳ1�>c��Q�S���ui)[��:�3�ir��A��7�\��j�H�k���s��RD(�v�7��j	#ht��vWZ,���i�8��C���ى{o�wn�9�՞u�u��s}�0���#~���Y���l��@�9��bf��H,�r���-�B3�r?�7\�����{1�?�M�ߦ9tݢ�����/M��Mjc�@�y�"[`uuuI��Z!w[�A*��)e�x�¢d�`di)ب�^z%XQ7�m֐o�3E�*nF�aBuad�m5�G��VٴD�):.Na\�*�R
^���������s���E��Y��Jq��LT��6��Nf@���vJ�*��b_��������I#����� ��|%hbT��.�����K[LF�矩%�k��eINd?�����k)���>���?\��3��XH���T9���Dr�;;ک7��%�����O�F�M�Aʀd.�ZN���_Z��NF4�`�1X�0��ɲ&!���\�%	ٿV�0C-F�e�ux-l�_��0�ק� �=��8K�T/��kzr��O��)�S��0E�ύ�z�<�ű�LA�P=��|g(����������"��ŷ'Sn�s��Id������=�"�V^��;�̿��\]+.����`�>��9�O�|ja�O0��+Pg�nP�.{:
Y 2�}��`$w�P��h��fW���d�����6Mmtn��?8�ۮ��U��x��(�)���5---.ۖ�8���2f�XJKQ��ϑ��y��G]�������'��,�����)��E:�j=~���Jז��+-m�]��������bA�b>a(F���raw�[E�D�e���߄��9�Q3Pn�o�دk;��Zm ����/���U��G��ueƴ���ܽo�Z�3!�-7��Q�q�ͺ�w��V��吇-[�����á�\�(՝r�Ţ�J0�s��|g!\A�Z1y2�7�Vtx���YMlO�;>��i�95�zQ�ppp8f������%���LL�ם��PB����g|--���i��A����H�U��� 2!�O�h|�5lΉzF���?uS���]N��b2BIP� ��&�L��o`iG���=2;kw|^�p0i�7`z16� cJ'jljZ��?����ۃ�������p�e|3�\9����t��L� ��C8��F���?Ϻ�Q�^�G3N���N�������wt*�Χ�T�zQ/''஋e{E[�R�����(��\MPJ@��Yͣ ?:`����u��iΝ�5��T������[xp�X�M	����vS���<��+�O)p�fx� �ߐ겊������Ҏb	���Õ�|�.=C�Z��7�+���B^�4�djt~��XK���Cώ��4t����\�Y�S�{⌋�\)��TfM�+_eҝ�C��\�v0�u�B(����ZY��F����
�ܗB-:z��B��)scӋ&U�d�ɛ34J��ۈ.�t��uc�W��gfO�mz�	*UO���Ζ���}z�V��w�ϧB�𱧪H�U�i��U�B�78�Ɉ�.;��?uW�}�H�`W�0�߷��q6�.l��Ų)�\���^Z1U�R$��6��USGW,�j�p�j�4����~��������}=u�ޚ���"bb?��?�,�Ժ�6�4#���������Y��ϛ�Ua_G�Г�LC4�n��������Sl�"86[n��ꑤ!�A P3��SEe���ݧEL��bc2�HG^^޵��#�b��l��i�=��5�3_9��/`�5?YNC���Ɇ�P��B�ľ�ee�;R}O-}n��E\D��"�?�w���f%
)��;�@kTU|�a$�@���%چ~�W�Gc���|n�ւQ����]�0��J�8ފ/��Ͱ��w�<��vW�4ͪ�����p����zʨr%YX��p��
�{�N�Yr"��͑����1�B��~F�f϶�?�O���l ���S*��:6���&�禧�a�wQ�)J0�n�m��g�d��<eWV��\:��Cͱ���w�6BxY�F3�a��f�K�(�i��v�ݼ��V[+�Q5��`N�ix��\=��ߠ��m�\����ҧ����=�(�S�(%R��}Դ�繖�t
��8�Q�eL��F��m���L��`�-����и�v�]��b�X*y#�BCCH�x���Y��44�B�|QY���w?����>������� @�F-�3�R����O����R��ZN�9O��Sm�s��Q�`� �	�-��ʽY��C�_ѵ�R������<��2�� �n��7v����ͪN�wxҵ����%��QE��.��	�֋#w�8�"�j*��5�Xf
ٱ|S=���q�����ߔ�~,)����yH�����AN�e���-�P?f�d;��7�����!A�f �B�Bp'85:���M��D�%U��|��N�"����K2^����z����� U!���^�����Ey7x�fW�G[j%�2�Je����$XP�"ԫ�ַ?��0�۲��^�`�j$�Z�9>Ģ��/��v�M�#)����C|�����O�m��»7~���1�ս5$�\y7��խ��YcB�)�e�F}� ��g�[�33s��9>��/�����/(�aggWbL|�D'���
���>˧��7����y�%	�H��*|Z�+���ʊ� s���Xb_UI��6��{��b����`�U=tu�ⷈ��vd���h�=#n�	�q]fE�$�W�ܳ��ބbG�*Yh�_��=|G"��Ǜ�}�>���xU�qX����B���s���v�B�c}�ҲS&6������Ď�Ȱ��@�@X,����*�����͜㻮%�=�JY|�UÓ��B��Xp�͏g<۝_���s��W�9O��yƉ���|iރ�EF���(�I)�� �B��b�(���{-����eW�dh2����"x��<
����dM��Z���>۸Z]ځ��.��e�ۖKY�~\|(K�Y�t"c��E�}8r8D%+�Dn�&zk���ё���/tކ+;;�=�Z�v���æN:`+�1#��� �d�IyS�i|i�����M�r�֝��T��>�T	�K� )k�X����f���u�&�5TQ{t0lCTo�=�A��e(��%����/J�J�\w5Α�t�Fs5����h��֦����"J��<���yVi���]���EHTF/@���ɽ��r�o�&+[�NP��u���/�m�lll`F6�G�/eP��
�J"""is�R�����˜n�\�����+7��!��"��C�qT���mL2Eq�nzK�k1�(մ��Z��0'&&�=;�>���#S�D�x��	*޺�#C�����Qh���Y�듛�{k�<�������Y�T��2�%�q'�+�n�/NTH(I��Cw|��"�
ϑ�sWC(��Yg��>��	��u��N@E���Ի�f��.��>U�(s��*�>C[��mi!�A�,�i�0����6ZP���eb����݋2� Į�Ͻ��w?���d��Gl��
��2(�P�>#�]2Em_~��M[A_�O���G�>Od��mm��X��fN��O� �q�*c۾>�u��]�6f�Y�[j�q�4���1��2��%~���緣��C��<�V�x[����e�.�J�d"޺V�d�j��lzV��E��{�(���%�6�w~�i�0��PZ�z��,��!���c�u���t��&�~6�ٗ|��2T��l�QRn)���\�T��c*%�&�-!�׵Y����I����;��g�sy��Eg���0.Ѽ�v�-?Κ��{��א�[��lCXG�cߥ[��"�2b`�à�J��v�	�u�Jp���
�*����O��^�7��^u�+4=r�����Y[����3�����w[D�N�"��/ɚ<v����(��8������0&o���{�2L�G�Ր�Ϟ�L�ӻ��p��o�.���P�l�隥��^�)�Mo�p�	�j��)��LUy ľ17Ρ�0O�+\� L�gQd�a���}�2��t�yJaX���v7ؿ�3J_����9�]'�>�|w����W��9�,/�F��9"'}۽+Q$� }�:�Rx���5��������c�x�Bw4p9+�/�
n�'�ǐ���𷅫��������``y=���E��r\X �1�Ɩ�3�Z׷�t�\<���y�w��қ���&F��j.���./KM��m��{��h@{����X�:��@���Mt-���z���ݪ�Q����F(A�>@�gZU�_������!��h��E0A�q
�5Jgk�_`�YJ0E��{F�8x$i�ƃ�d��ݨ_��|�]ן`ȗh��B�r�}�<JSn`�5φ8�-�ن�A���}��� ���D�d.FW�M&�_���=%^��0�R�)��44���￱�h���\��CLJz�.fdn�ޛA- �VT����1�Z�漁��� �i�E�4R��o$���E��6�Q=ʂ"eQ���^�P�����ԻJYC�s��)��(�W}!:�O5	�޶��5|�_4�<�<�K���ܩ�;��uus[n���Yw6U��EuYr2�}�L�Z�o+*��N�n5�{" �+�B�G��ۗ�T�c���{���^V�ɕ(���w�LZou���SW��\xJ
���f���>��hhh�{��������a�W�e��0\�M09o�^	FF$IXɠ��fo����� ��[?���t�k!􄲋J�Æ��P3��u�;�}�W=e�%Q���T��G�_�b�	�5��;eD�$r�,V\>n4~r��J�����N���k��ry�3^yU۱��-M������_�"^�'1�}mm‧�j�809~�P������xCq](�y4����p����my>\H�ŧvKݩhv���������.a�闵F����_D�oW%p�&������~�x��g{.'������쟸~&�ny�Ē�5T�֎Rڢ<��gBj�#]5��2�A�BbF�� ��7��G1.2L�Ȃ�%��9��-O�����7e�i��A=j���\��A���Ǜߑ��Ǐ���0�}S�8(/jѦ6�m���P���v�T_m���[��xxŲ\B�[?�V�s�����G����;vr+>� ��,��|p��A��[-Sq��~�e�U��N93�_���uUי�x~~�y��H�n�޲�2˼ʙ�r���8�0'{b����2��<������lH`��ī����=�5��E�5���A���N�^�[eN(�&�t�1�)Wӯb�.1�)Ƃ%$j��k�6��SMc[[���b���������^�`��3Ԑ,N��e.ҟ�y�2�}ޣ���N�l��f��6>�Rpc��4z���Tb6��-��v!�2��f&4�ٓ��U���"@(OrGN7�ܩhږb���lii1�fd`Px��zl�������2�D���	U����@��g_��̟��?��uͧm��E[W�o;=9-Woa�������H� $��,P���0⧣����'���cB8tˬ�p�}�у��^�|9)��2��EP��DĻ֪@uB-FÃ&�<�&�:z�n�z.�ީ.�>�Y�~�ܽZ�
���w(|�#H���'�k������fE�:J����z�CY���uܝ%ᶬ��x9fh���Z�n`E�S&lE;�=����;}u��Rm�����e��*��7qGB�|�(�����}�/�N�~G��V����?�ى{zz����OT5[ES[���s�\R0\a�X"�Ng�ay0Q� ��O�h�Xn�Y�{�e�Xn�48����ZFD�}����]�W�TܔG'�j�k*"���>���bۻ����f����4�깔6��|���L��vN*����M�?�T�J��lZ�fp��ex����O����R��R���d!�_�7ir_
^�}3���t��ฝ�ϐ��8�Eы���W��2�D�b�yy ����4
qV�.-�w��Z�N���U���O�Dޤ�Y�/����3��Ȓ��L\��.�W�xbd4P�� ������s^a�u���G�A�d�0�ŷ�߶ܩ9c4үe�Y oN�Wd�(�]����h� T u �s�s�#�O��_&��u���\ĥ����5�
&	�ϖc����	����#�j/�⌁L��cj�t��܇.٩���P,����Sb�� ��ǐd@�w>]2\c�Q�Pz��Jf&����9B�X�,d���#/}��'�ꍑ���T�2�U�����]"�l���dP�����_�nV�3K���������ϟƻ��!-�F���^��R�J�Gy�uTD�C,@~{�\�~LT3�^P����t���My(t��u�(�M]Q��X���"k�����~�����F֖<j`ڵR�x[���ן��_h�ɲ��)a��[jS�ѿ��Լz�_�����W`![��C�BB	G��=8�����u� ����R\�Պb�U���[\�Aޫ}�`Z�q�6��,�<u�W��q�0 rx��O����T-�e�yN� xT�}}���}���8(})S� Е��e�t�YB��j�U퐎Ŭ\���`0=�d{� ͵5��Z|nVba!���宐��F�k�Xt���{�v��/4�1��?�ܑغ�.�xp˥o��i���s��X;ѣ�'T�5;%�p�@ÜkvГh��ԁ�˺'EMWo+!� �ȝ�vdm���>rfKY*[,9&W UZ
<%�~E��N��G+7�y�Q�qƮj����{YC�F�ɔ����}�p���Sn���O��U�p�<Ϋ�?���IB t�/؅��]]tU���l�|�Y؍`��'z8�l�9��*iHz��| �8��Cf��ZH1����gWь�7D��߿���|aaa�-\�>�Q(%5>�j���~Áv ���,� �q,;�1�:����=�z0{lcgו������(�<�bQ�}>n�Wh����NOg����6�D��*������9;ϭ?v��^����}$��L�D��=1ߟ�]r�����qj�+]��75Y����߀��-�Q���۾~毞s��S�1���0�J, �3ӣV��I milū:�o-�5��0��v :��3�2�K��u��_�������]W���Bi�z��/onn�lR�D/��
�L��Ngj�?8����ӊ'0���֯?���6dD��9��.��evD�t<������2c\���^N�u������_�Vd�������gZ:w�,7ch�M}��� 3�'�z�B�K��o��tqj�c�N�Ne"b⡄g2�ܑ4����^�����4#���k�u�v�O˥�O�+-��v4��;�Z��'��n+��K�(��_ރ�ŗ���ҷ�����R9�GY�B���`��D���GP���TEt�����e����l�+��@a���*���.uS��^�R٨t��3������|L�:m�9"�o�t�;���>w�V�������	d����sAT)�������_�x`��XF�R��,�F7^��7�+��0�Ҷ+��>x]����$v_)�U�(�Z{/*ޅ�LHF�oe0r�}�VO��L��H��m>��R�'�F��}��-�j:��~%=$S�F[�F���T_�Ɍu~���� V4꥓X������L�E�Q��:�Ζ�ɼ�KP�t]��M	O.`�999A�*�48CV$='%��C$��߿�Js�h�`� �R�R�C�V�S��LŏF|������N%<`����� ]6ֈ#KV22���u5�+7h���G�4�¬4�������ˋ��.&��Ђ騟��.3­�J[r��"R���z��B�����J����M�	=�o잝�D�\C�*
(e���^ԍ� �7X~J�Y��ELLNfl�����"��Á�4;Y6in�F�) r�qV�zV�m����_���j�1Rb0�N3AW�D�;@ݡ��_��~���+o|Ž�v~,	���js���|�W������'���Gd�ם#�,N�5~��"���<ɏ�����C>2��������A}}j����I��,:Ҽ9�����Ze@[&}8��kv�H��$�WfWx2�~�@K�u�m�|�.ي��@�:������04*�w<�k9?���Γ#�g�g��� 93Q��E6r 	��|�Ao22���]#~�RD��	gs����oy����p[_���<�w(�M��Z*Eܧڼnﺳ�HL�Y[q�9�/�M.����Q�^�,���E�&ƭ9(&&&�(�zEr�A�3w6w#��͍{������ R�����X��(l^E����o5��	���x�v����(dmw�d[�Z�6C��Q�׬���F^[_��1^}O�;����m��&VP�?�|g�[�{��$�q�P� *�֟�yFf������4���̌ #����������#Y�
������Fݗ�4"���}�M��o0���S&����Y�V�＆ګ�6t�����FD�c@�-j�kgg7]�*����+j����/io^�nʡ8�J0�1���m�������*k�ֽ
�L�����^؃�k�b�^,�B��ONҼb�e`���U����	����(���Eˏ]�����o(�F��7�H��+OS$��I��|T��ֈ���۩3K��Z�����I��X/i}+V�"����J����c�<��{��ؼ����>�ɨ�yYl-��m�Tu�?I.Ds�#�y���H�6E>u�� ���	Μ����D@�xCCC�jZ�sN�H���^�ϫF��M&Q(�YMMM�3źY�VHjQ��qx�[?���w?��T S�B��e��?;n!i��g����|���ů{�v�A��&S�j	�R��/Eg�����!ׂ{�h{))���mC�ߥ"�޹Q�f����0�%�CU����*�!���?�����E�0��45|�3��IJs$�l��s]��b�C��ÅI�Q5�[��?4�8�p�nE ��_�W�!)Vn�@Q�z��Ow�<&A����h.���ܕ��	�u@D�$�;�l�b�/?��g-��,7���S0W�>�� Q��=gK�p5Y��Б�������oj�v�WJJtnO�\cR��n�� �թC�e���t\N�_jܨ�����Βh?���:ktۀ���d3"�(����l�+�	�Ό����'�3mx��o��TJ�y�",�o H���1+��N)p��
}W(�Z(]��ېВ����0��@|���n3h�e���=*�1�O-̴�ٵ�ˠ��z
�I$T���zRd��RP�cz:�
�r�F�0�@9���?�漊�~R��PVk�K>��Ao�r�w�P/@�'�I�Lʳf�$��v�'c��дi!�y�(��Y˔�6V@-��ƮF����-�ٓ�T�>�^ QS�.���zYN�888��a ������yآk�ǫ��Z	f�	%m�ī�PDP�jJP7V�'��c��J��0��{?����v�o����j�r�I�4jϓ�֭[�jP"�2B���H���[�P���고�W��}#
�+���gw�~_�C�8�%��hvn.Hx��ԝ�9�?�i��}-~pn]U�����X �{xH�O�ɘ�S��e�|��Ņ����d�A���Ž�m����-��(-�Z���6��^�¼����#sf���D��O�ـ�K~ͫ��'�0�tE�b�V�p�a�,�ZKb(وn��C	����b(
��߀�X�b>��M.���Elsss,�)U~*��xM�)�W��Ӄ��U�<�AO�q�Ƌ�B��=���z��H~��/:��T��2�X)o�ÒJڲ�s�w��Q��>;�็�*����$x�n��^%A��]�g�J�� ��I=��{WKMǢ�rƾ�4�Xj~X�JE��?88�z�S\O��S�ea1�P>��=����=݆�)ѥ����!�	�&�\2ׯ��.��Ȃ��Z*��_F_l����R�^�Vrw��T�x��P:Q�(��ׯ?�ǖ'ÅN.������t��j��HSSs�3�֮w����v1y�2�:���QkN�^5 �z�,�^{G1p���:�	�s��p�V�z��}��f���Jj ����x�����0��/ۍ����S&�[���cK�Ov=e&x����v)7,�%�?2�\�Zf�'�g��Ҕan�|��l�����8E��#v����ͱ�n��4�r����p�J��e�R�+�,%$2L�����]�a��b�t�D�� �{s
+=[^(��7/E�Fq��&�̮&@�զ̈́�Fz��PW7/����\ V���?�1D��J�9XYAg�����KO��fB�>�T��]ξiK�0��"<��������=;>6p3��|/�G�P�Ku6Sf{f���&=�~d\K�ƙ�0���E�(����E�k�?ᛜ��+�����;G��`�U����N�5~_P�Z�m���}==��ʾ��RS[{)F|���<Wb;�AN�v�YW�m��kW+�X�?�,�k�Hz�H}5!$�������f��ܕ%ᶢ����F���[P>�oM�+�Ʋ�Ȕ*�jd�8��<������j�fĠ{!�/.v.� n#[�a^��&�/���)�	�H{{;z�5荬�!��o�udۧ�� ѢW���7�⋓oƿ�����/GG-�-f�ر�,2�[�d,���$X�D�Oˮ+�)sz�fr`��m�w�u�l���1>C������"�H��z7P`�ﶻԧ�]�
�����9F��z��l����lJj�b��&������(o����Xu�?�l�N��r�~��LNZn��'��Q)<~���%�CM'��C`'����=3?~Tu؁�;��q�,�od� �xE[��m�^��?'y��@
Gp��8j�U*�!�Cl�k`1����sqT砘�t��9:��/�imc�#]�В:&.��۱i��2L��**��B���+���&�P\��fc ���5z�y#�����4�ty�ْ̆�g�PG����_}�k[[uvx--�Pi����>h	�/_�_�PM���=7'����G߲ZEe,)ѳb���y@�3��I
d�Uv����%��v�{oB5��<���'{?7:��x��iN��&�VN��*�f�P˨�}V��N�ZT���{]b|�߿�O���1� �؞m����S�Zh,$~Vۼ��Δۇ�%A	�Sn��g��ݚfr^o�h ,���ۖ���	W"��x���J%A7�jx�g�C�)�JÅ7�_%�a�Ky�-V����1������u�.A����e������f`9h`9��D�hc�w8JD�?fg ɤ���;�ޤ�2�s��U����N�΢N��?�'`9�7�8::Nb�.�mg�v����wL���Mv")|��e3z�Z���~�,�P�Vj��}�V�ƕ����%���̧���Fi�ؠ�д6>�F��(;D��YzT����h1e�mݷ~�[Ѐ/�S&G��(~�*��m��С�-]��t�l\:I�g���5��5��q��(�k�0�ž���HT{���a����p7L��eSn����a\��GAr�S-#�v` �}e���x��϶���A�A,/��x�2*�@�e�� ����O��x[�P��8
y]�H,׺~FK6 �nhh��Ŋ]��-:zz��am~��k��^A,T�P8h�DF���L�$;f9�A\���_`��>�[X(�H�f��������<��fٗ�yu����"��tI/ � ��YHѶ��a�q�����r�4�]V��D	��N7�Ǧ�e�xY�=�u�=�5�F%8]H��k�И�5T���������T��˩V�Ԙ	��7���G�H��̒r�9;;�<�-��8�d����#���t��A��%�%fjC�'VbZ��Pzz+�������xq��5��u�@}{Ɍ�����l�bL��;Z�ߴl��.k[���9�~���Ǟ�����ӧOWs �Q~[3�Cȶ��ҵ߿��2KIKC(v�6\�y?����/�8z��
�Y�����YPD���$�(yK#���;�~q�s�� �o�L�~� ��&�At��t��p�;��� ��EE����@�Kژ��5V�A�2�� ���^�,:�se���Γ���X��>\��@˛�!7������ff�r�qTF��@�e�q���&:�y�?ll�����ŏs�8ɮ�<���4ǫ�@	��I�+]�2ï�	YQ��QMPf�vi�s*���wParQ�D�6���������/����8_��y���HLO���F��^��E���^��~^��T^-���8 �|?�����l2v��)�d����=.�#%2����N�7��V���^(]����`%-xm����X��( �K	���u�Le�(�9]F-o�d��o�R�}ʀ�i��$����:�n����u�P zKKS,�i	x����nz��^���lO�Y�A%VtιT�X�Td�Q X6�Z�B�M��銡�U!���=)Tǫ�|%��<v ֋�s7h�W�e.�E������v����딍�e�^5�\F3����
3?��j�w=//��=7YD58��Ă�� �y�w�t�J?).�.?cz�t�z"���6�iK�\-�~�&W�",I�F��g+�dn�������<R��7붦����Z�bP4bK/����m��_���%�d{.�j�������[��w�,��@�c~�ը�-��B֧$a�c��C/N�f\��j2�h�\��?�[�t�2Z���n~! ��m>p�$�*a�����6Ƴí�yk3:@���ϕ�˲���9��ΖJ�w�����=�
t�����|��C�!�.�}��g��U)T��^u,���P�𫥈�ee��ۉ��=e��f#������^���bĢF1绯�a|=�������C�� Y�B����~||�d!�>sm�tj?��% 4p�׽�]\�q�B�&�Q�L��킧P�)e�2Y��U�mm04���+"��l�VY�)�h\��_W����I|��ʺ�>!��ߛ��o=��+��PE�����`Ȃ��?����r���EV]]��r��o��V��Ž�|�\�_�BD��*����ޚJ�{�O������J"�z�򴼝Y@�@{c$NE-��UX*�Ѓ �;f�8��d~
����"9�'�Reɯ<n|6$Ȍ�N߶������1�̤���!ψ�������)j_�-�?�-�l�H��UM��ppp$|��^� 0��9G�xGa�ez���#���DD�u3�(��,*����ؐ�;uE���*Y�;�/N�I�ڋ�<��w/|8�*���g�����X��(�a�3��lv喖~,+�*�1B�o�$�:C,yq��[CP6��P�F������|�����ՙ.��/"H��l�m0AEto�_R��}x���U2ݼ�ȧUB�h��㳥�x�CP*$ZBYxV	�x��2�>��p�ja�`y�_���&�o3�	���9sq`'�'@)��9"��)������{��L��V�:�m�٬}IO�%��7�AYf_�mď�3��x���H�*[/dZ�8$3*+�����N� �T���{���-�n�/A����/n��\I��F7f�xv"x�ԛ�W���P�Cz<;�v��ni�f;�Q$-����I���f5��(fvv�;8-)��"G:{��tM�c�1<v(���痏.i��!3[EB��/\Mz�l;���ۢ�6���/��ý8���Z�v�E�Z����ۡq㮌e��N��r�-���FFQ�1�pN*��|�xUJNF< ��8��(T{�W.t�u�����
���%��,�g�tM3W׉�3���4����N��fW��&@��yHC���¨�WǢ��[ﶢ������ ���#M)<��@�5a�.~,!灑���}W����N�v�P-�
N�*.�g�w#����8����r�y�^���#��oWȑ�7zZ}8�?��n<;^xў:���Xؕ�!(�k�;��V>�0�Q+J(c�iX��}qq��qy�D��,`sG�ĭ$���*�SI� |wf��0y���i9ZZ��[g����u������ytK�p�` �Wk����"����<ɀ:>42���[~���<{�z�/�3�h��d�wy�tEؼ�����c�KKźD�&�￵7���}I.��\1��א�$\����z�5�[���}I�m����2�����ۊ��A�ug�6���� � 1Wz]�Wײ3ԗ�x$L.��^�%8�h�3���i ��XB:@W����bbb/;���ԩ6Itu�=��Xi�w��g4_�M��y��#�������~d�n������cI_�������}���IX�m�~e(� t���{���Ts�aZ���8���		t>��^3��#Sww�������0 UJ-�!�}��׍�ЅE�a斍���M�,��WG}H�!տ��h1�W�o��m��s�M�2�I�߱8�ߩF�s��J�����i��P�,y�o���8XP��d�!�8��q@�h�c�˽�q��-r	g����Y���9�0����=Y�o�u�QBSài�ܚ�Q�Ȅv�z��{�+�:�h+��	F�\c�/� ����#^)3���P�/�y�Ih|��kG�moo���}������f&��~�����sP.���e\�_���ի0����׽��خn��J%��KO�K_8%cLmneYYG���`��* :O�:[py������n�A�
R��;�>?.�=�-;iǦٵ���H��ܔ	�P,�g�����~z�z�vC����Prz��Ol2Ū1�� �,N V��)�j��+��A��޾J蝱o"�c9�����A65�5��)��;455����Fc��&�s���C�{��S�w,��aWN��єۂM �y_�y�E�M�gL[CZ�O�5�8����މ���]��@�]Hs�m7��]TF��x�9z~z ��:>����J��6o_��E��2I��z��#��Sy�ұ�&��������)	%�ܛ�T�l����PTѹ�mX��R	"R�_����V6�M���	e� ��(/�T���7�/�%�'�po���h���d�I	Xk��L� �'K&�r�s��6Ubf���.9��������>�m��\�����`oMtWuAQQ��!�~2��?�잻�x{c�����d���0��Ҳ��� ��Wj�V���g̹ڌ�]�Q#��2k�*=�Zu��VVV�Mmd�zhh>���v�� ;&'�����8�t��r����u?&��7ocI%��������+��xo�ώ
лi�g�7q�g�ɓ�B��i�	�`���bg"#o������X��O��gQ�V>����Ο|������VTV6��^p+ V�^��@�ul�o�Xy���� CB�#3 W�w�B4u���Z���q4�p��$�A/:��� �0�o���� ~��5W~c~���<P��Nfv�&U�ׯa�&S�9.�J����YVl���=h[ށ�S3�Kx��ȓ)A5E�3�SzQS;�ؖ�W��$&u/�C�����@�w#���&��$a+������{�cV\J2�l
���[B	�5y��|0ixI��i���U�n(��TÃ�&��n��V�E@4��8�v�[��lH��v����x���η2BŜ-��'&'S|���锕��KI=��P���`��C8���M��8�{4,
�2�]~�+V&���l�s����~s��wש��|K%�k�C�)�����F�QހX�ʊ%��e>���E���$�R:�뿺���_�8���t�"�Q�� 짨�a����?e��r*
�GP�0��v񭌢��������D�F�!�rP}h� z�za�!�$���!Q��f7o"P0�6���n�ʕ�2.�f�q&�T/�7*ۘv|�Ϫ^/u~�v��ӻ��Po�z$}�6x4�%�µ��}K��� ����U�vB��&.|�WWee	�یC�ǹBn�m��7r��Z�݈��ԪPƧ�M��R�C�Ļ�Hn,����o���+������2y�������0hr��&���������������y�FZ������U�XLB�%�QR��EbiiY%\���%TD@$�F�A��o���|�=���>3w\�u��3ϯ�ms������ș7$�����6m�أ���_���8�e!��[�(\R����� 8;:���?���j7˙�|�'_�xhc��;\��i�;5� ��Gך��6eK�C����Ӵ����l��!�2�>�u��_`g��{:�T�.��#݉T��?+���UK�y1F�����9�j��6��̸ W�^�pƦ(Z��NI�X���!?�"Qb>�su}u}��kM���k��,���=���9
����7�L�ݽS$x���� �J33�u�s7��(�QX;�fP�7�ػn�'�_��`�	�\��E�.y7,?��t��5����(���=��!/�nh�:���V+.>#����m`5�3Rܳ	^K���]�9R�bee-q�V�nTϼ������{*.���}��3��"�WpL�bV ��q�F$
�5�iBd�u���"��/���ꆾ��v	_kQ���Oo'>D�y��9�X�/bFG�&��)=N���~�����u�-�͵�Q�hN�c-�U/bŠ8����[7���⎦)�qQ�_�C"�4<0ħ�8�����[����_���KƟu�6���e���d��(�����nPC{��� fq}=���/�{L�����j��&�C+����0��D�h���X`�rU[�;%K��~�Y��G�mx3׶G�~`��Q9Q<Vg-w��$���&H��u:u��h�5 &é���+�ۍc��kl�Y4G�"Q��G����)!P7���F'��ӝ��������'I�b�@E�"�d���}敢s52=L���W����mEM�*}t������c�rB�7C+��?�؏�!��}}}�G�����D�ء~(M�w���gE-�@�ytbNEdq�s+���K������nN\�o�t����4��B�}�F����w{�g(�
�{�G=3*����xM���C�]�����W*ؔ�ۜ3�#���N�O��8��&[f�d��8�6w��^Uh��~yy�9,���ף,�lS�;��/�� V6�9��n�F_@�]W���9Ei��8��4��H�����WA�� ""�U�`��F�h;T3tݐ[��}Z����\��ƞ�'u���<��۷ob
��S�Ȟ��ܥ��u���j���*�ٔ�3����ܴK�d�V�	���Z��*�Q����`�`	"�|pU���?�:WV&0��2ΐ��^H:9��wlQby˳Ĭ�P��9g��]'���B���AkJ��b���ۉ�U�B��dO�cN�[ݻYu��ne�?ee]����t-j��ښ����ʟk��1���+���DrU6�`|ϴ�oy�(9���%FYQ]s0��瞴}�[�egO̬K��Q]�L��:����:�A�5[�=S�uޛ�+��5���k_�/�@�0���L-���X�Q��*�e��5s��ӭ����qݯ�|�o<ײ�}����(
��;e�f��VIlU�9�\E%l�Ut�l���c������px��ghH�A�#��?�M|+�#.��7�JWُ۬�qh��^����uզ=���f��m��bɃA>��7x��S��kɪnI�xv��/?O�9��Et�_@�4��YZ�u}���-2�Ň�=I�`F=6MῙ���OW 5��$�BD���@�h,t�אD��L�Ũ�)Ĕ;Y��.��rĕ���
F��=s��^ �����p����ѽ��_˽i%�H�u�2b��q�
�p���뤼�����1�rm��|��їDj���3��y*�5|]�vʽ�J����c�p���������$%NT�NO|zk�B1���\�����&.9��1��B��������)����I/�>��|x�;��)��}���Yh��CKP��Qg������Z���(h���$��٧v�$<�l �L�V���?+L�K���!W�a{*xe��|&�x`Q�\G
]-n�_5�X�IRe�>�ȕ!\�#�]��D��弟���:he��Iб9�Pkjv�-�'���GY-���:3��͕�Ks.FN�l�������(�Я�����	���Qbr�!�ژu�,V�NSUL�Zd/2�+y5$�:R�[���۳���I?f/��*Z�S��^NɁ�� �`2�{������	���>S���+��#�g�m�B����7�����O��h�/Xf��6q�I�#Df�i0k�^xz2�YU�����͛h�8��d�����y�����sO8/4�\�E͋��#�/�qN�ErY���G���rR(�b5��Q@n�������u>d��䆎Rtww���u[�z���9�c�l7�wzzV�]y���JJD`�ij��R���r.D�����a娰�� ��E��O�k����P�k@�vjy
�ze��z!���x/�]���uDD�C���a�AP��`����߿o�?�R扽�M+�����:�Z\L,�SFn�Ewn����˕���Cfw.�:�T��X�UG�j����L6�S���I���w�u
X�~4��^b��/�93�/j|�:g��_~��1(�f��{��U�
��>ܴ�����C�D�.qƐ�]�N;��`�Vf`�d�����~J�Vp����d��h^�[�fv�{s�8�W�0N��ۄC��b&��p(��0���L�}���U�#���Ћn5��G��0_�}�a�[���M�^8wJ=�ڼ'_�-\�?�&-]�W׮��ၼ�=u_��9V�.4������6:u���d�W�ݧ%.x^I��hת��>��يk�U�\����U.Wk��~u�m'�7�7~��h�0<�D����P��h�q2('/��T����%N�����c����S=���v[������y��K�r}p�g{~�M2(��☧�N1Wfxa'���2��.Au��s�Rf�Q�e�=BCGG"X�*FD8`�ܒ��P
�.%��~�_�Xk�}�U8Sc.=��j����6on:��}d�&���[�9�~vJ��[�VH�����P�7��t׌{ص��Z�M��l>e
٪|��Bg��;�T�M�G��zHc�L�Q��خ����C��G{�YJ��'��)��
����;�f�G�������?���on����^�z1��Z��G��cub>O~�����r[}�!�$s���6
~n.�n刭#�HE�1M��ٚz�bs��EӖ�W ��M�����/�G���)���be[����0+^����Z�!�B�%���s��Wv����b��/_�����<I[cw��Ů�	�Ŭ��X�Й��A�;�7Xi\;OC=�8��򞟏��x*���=�[�o�;��Xr5��(5�!����΁�._����VW)�A?�j�'�ק�	S4[���%��;�%-}ֽ�)#9y�qP�Ҵ?G�k�.|��;O�������1�)ֵE�>}z1V'.��Ό�Έ~������2�Z /6�l��������dx��e֡���_�u?5@6�+]���HA��w�?�jc3�d�RnV��,`��M�8\W�<�L K��L���^���S�W)���t���@|��I��x��8�ӿ��>S���Bfouy0�|�iC��kZ��ţ�����,�w���w�\S}�b��?.s�?��UIz�c͇LL�	3C�^����-���pn�ta�ќ���P舃�߱$t�b��������h����������g;�t�^~W��z>�.�@��~d��3c�C��VGj�{Nf$��<)�z�nϕA�=mo%�O�Ha9�d�^V�N��G�8^ȒX�/��7,~���$&^����N��1@��ǻ`x�,,�K�}��$P�ȎcȞ��+#)�|�pu(����ג��B��}cc���?���7��w�6��)?XCh��ϳx��:�}w�j4��p2��C=+<�ַ��Jr���L;cA\��J?�Njp����@�Yi7�}:9q��DtF���[���'�ok�IW�%}}���Q�����rP����ōg_ X:-���q����b��Ђ�G|�&|2dd�TX��1Vɵ'��<,; Nm�Ψ�}���DI��觚����QgϽ��5�����z����@;���H��0t
���ts||�V��� ��"�UE4����}���'�R�y�)����������ټ�w5���������/1�r������.= z$ ��f�Q�B0���k
���<9PM�4��J��鄙�ڭ�����od��YV��9��J F�(��U����R�?��LV�Y�B첨�O��o��C�7o���QRS����}��]����*���⸐R��K��ED`p��F0�7\�T9�Kf�L�#�|���_zY쎹;������N����Ԫ���k�E�{��1��uΠ�?�b~�����gD��ǫǇ9�r~�![�vUU�;Ȓ��/�̤e#׷|���, �;x���ć ��	�q�0mL',���%�pyej:��	���KH@|�ƍ@���ﲈt��rN��}ХuĄ��y��[�IZ���R�ҝ8��v���/<hrKO}��#'>D�E[a�[Xߚ���R?���1��{37��o��H��]�{a�IIL����B����5����k	�`���2��R��B�8�3��M���Ukɕu˓�ϊ�Y�[�ܑd�'��0�P�;ZB�>rƔ��_����4@��l��,x|5e�\t��v��@ �������9��ee7c�Cל�׉p�%�B[.�7mɀ�}��ة�rRn����g|O����W��5t2W���7��|f������l ��<M�]�s�������k�#�~n�����z�C���y���GT�o��l��QP���nCC�Y��d۶5	�+Ýdq���>�E����|<�X�j���x,�[J6g�Ώ�^.�M��}�� �t�C_����@;2���((��M�#���J::L�-&z�u�)���xQ����:qEX��9F�,�q~�2 DS����g�	㐗��>����Vn+��zǑ+9�8�6@���WD!�c0[t����-%�{u%��J�dty9=��1y�~���Ͱ}�s�x��-S_�AQ�
����M%�����P&����b�;�V�'fZɊ�ì�;~Eo�)d?�����	oʝ@n���z"���卉���a�	"��Q���������&�gu@�<D''��VVj�~���t2�B��=,��� :�jv��n�hI�X9^�}�Z����!�{	M�W��l����g�xxH�^��P��B	!h4C��l�o��L��[��V�G-� ���U�'wLǚDM\���ؠJ��Kʴ��\ f�����4
�0ď6�N�C�ʓ"O�Aؠ��ո�T	t2�#:-d�`8���R��{��"I�Sp_�f̤�Y��ddv���"?��[������_/�|�B_�m�����'w��)J��P9d�����s��>Nkl{K�.)��u��@�a� ��F���T	CQ%%�_��v�)��k;66��8�D!�k��9�H��T����D�"��2���4��z�0���*��[�LeJ�����5�a��8)f��.K�Y{KfR���|�<2�1�u�s��n�/��Q���HD�H�B�3HeE��5]��?�?�O�9y��[�WOկ���VM���v��S�7�O�Iٙ�99:�6 �w	F�R�`�34�]rMl(.Z!'}]�)�|�� Q	��j�rs�|}}�Y����J�gP�F�f˥T��z�����[N#�J��'lg;R�K�dxx�!�Y���� HT�`c ��Aѭ�������^���H���(���f���eu�â�PTW�)�[��eܰ}�����Sr,`ET�te8�z於��4LU�Q
<q+�L���D���`���L��au��io�%�eDy��E���y �i�~�K�Y��z��e����x3����픣�S2e�������NM��{�%˝�p�c]��&�r��5��R'�>g��U{g˪l�O��{�7���۴+a7�{.�W�������� 3x���g-|*hbe�?�B�w}�ˮ2�*F�VZr�զ��KC8)�������vkOZ� 	�?��5�����OB��40�Yu��/ڭP,�����$�n��βc���'O�
���g��l/�̝�P�
���ǻ�
��q�0�=����<722�;�+�h?��E��iB�G{鋗�e�aݔ��&�em�ƹ�6<qR����������W�X�Е�1rB�{�-�7� 1���t��8�+��@��Q ����sE��t�픜+��1G�snK��un=0��B�� �%�����%�+mV����}�g?+��i=��)˛k��GZX��u�w�|�{R��D�z +7�qT��U`�PZ�r�����5��#�]��#9���-יK�d�g���?�1�
�'��2�U��j�iw7�E�3� �q�S$Vlj��.34oP�kY���Q 蹱�6�J�Ó���@�ؑ����ޥM�/��K��޿.<5s�rC�D�B�S
y���1Q��y��Vw��޳<P�%���� �Xna���E�bKR �?f��Q�9E$�qVnn(�0����4(Ea[� �0gn��K@]b�Xz��� �9!����,ȑ4L�ZI��.���ك�8�d�ȿ#��:s��~�t��6�������>YR�y���b�)�L��"+�Pl��h��e{q��7�M��n�jq9��B�:W�Ԟ:͈!���Md:ʢRy-�l7���$��*/兿�W�-�JK>,G�g�9��@�	�Z15ܬ�C!Fx�y\��\�ס9�;�ͩC�*Hw�my��J�^
	3M���j�9�i�=��>��u:_�m�u�c�3�LwJa:�qc�$�/���8��n&�Kw15�7%����X�-Cn������(# ߚk/6wt�g	R��$�[�W�L�;�/���g_W�lM�S΄-`��x0��?@��t���jz�g��nV_t�d򦾯o����Pډ�&w�J��jxg>�~;�8
��طL>�k�
ONN���}�hh��K�ZxeQ���w�-B�by�.��q��.6�J6>�(MW|�W�&��l/_�sm7DD�.;uO��)ٵWb��|x��C`�A��7ZP��6�05���|�	���K:Oӈ탫~+3`,�E��Nۍ����T׶Վs?ml\=���~�D6*)�Bل�48u�����Pc	�2qf�κs�fO��m�-޹��tȓ�ղ�����zeX8��B[I�IP�ɟ���q���Q�<�v���$��6Gjׅ�<�Ɓ�l9�vRL�ƥ�dO�(��_���j�����W.��U7xѣ-:�<)��j�\GGu��N&�h������oC處�Z�A��}�<�͑$���Y�>W|{yi�������>�L[Z����S*�*�J����k��X�V5sq'����J��� F�
$�<q��Ԡw���Y�-V��Ds��!9�����#�C��!z8�x�w}jN�����z��(�<��fVV䠐1VJz;Ÿ��!����?nbJ��5I�bo�|ݷb�@hCi,{kTS������M�D�2�f7ݫ��>I�F�$�e��w�j�y��
-�2���_4Q��oh(PP4p7XC.<���nEb
j�U��#ث��7��ˇw \Y<c']��ʻ���9��B�کo+{ͬ:���Է�A�fu��<�'�a��zEy��YKF��.4MҨ�cj�8�v%���><<|�2�J��ޕYh!������f�N���!+��0��Ŷ�I�)i�Y�]ر���y_�(�)���|`F�u��Lw�z��V�ꍼ�,�dn�HF ������S��
�%��	F� �6��@�� ����/(�҄f�E]�a��E�)�����`��-�0��$�2A�Q�A���u0&�B0���X�|�m�@G��_�o2�{���J����4F-�|f6���{(��k�tL �������̔���M�_�pjWЫ~|�}3,-�]	aqc���?=g�$��=*��_�_}��/2F/\FO~�P�H�m��9ֶqTyW������ì���ue��b8t���ڞ5�h�3y(�CZ�X$�;�@S�ҵ�����>D�������$Rְm2�u k�ܡ�߉X۟����rk�g��+e��:�{���(��+<)�+Y?�Ƿ�zG�"��H����,�R7M: v��wi�d�i��O�v��Vx��l�����ſ-t:��R ���3az뎦k��^s�������_
8���}2��;��!����
U*��=���$A��]�a��5l��T���W�|~_K�`8#�`.�����E���@�z&��������C^!��Ti��]K��,h��C�.!멠������I.�(��@y��@�
���5%���=��(���ږ�S6���=�ޒwxL�02�/:�JQe�tNd ��aԡ���r~Չr�	���.�º/ ��<:a�Q 9��^w��v�n\	�j\��Ȭ�N깻�g�x'w+%zh��-���G)-L�̨
���ٮ�2�[��D�#�G������G��.s
f���;__�3��U���:A�Mv���U�5
)��PW�1+�E�+kL�L��e	���h�Ccg����f�Q��~�ÿ�;�b�]R�Md���J[fVL4;^2,k<�2b$��)]q�5��黬�ǌ����+���䄼�����b��3�� �'u1E�B{Ԟ(`T7U�����xïL2]�S�3�C:%�ٚ�����'3�1��#�S]�O|��{�.c��S!X��q�Kz����-��9��$*�	���E�ՠ�YU�S�r�Y@�Z����k���㈑H�T���V�x�IW�J����2�(q�^?<kJIM����_c�L����s���.�Fa?�orR~���$��Լ��ҐH�kΩ�b�������0��E��}�����F	�Ǜ����.��ﮧ9z��
�q�����q ���1a���L��=<:���{3=mJ���'�B�� }WWWnfJ�SA-�~���� ��ǝ��aHhW�f�� ܿ^�����U=;��ïŬ :��L� 5d["�j����J����,��+��ke��¾ifъ�*=gL�z\�%���f1{6���)���}����-#�����@X0��}�{��i>�L�~u���. ���Ӌ�ט�i��;�F�^�w/N����>��\���@�q.��G���'	��u���v���.Rw|75*h�K���-���#��E��(���
�`��� qwP��,�pk"��T`�P��2Ӆ!���d�����$JOO������^��ا~s��5鑁��\,m��������F2޶��w�tۼ
��fYy�	�zI����o������=Cex0`׻@���m����"S�VT�~�B� TS�?�C�x�5tt��Q��G���>�(	R/��^	E�_?=�I�/ܡa�vط�b!�\n�+��B�'%
�����߷�0�}3x�� �[�@M�"˓��6�>���߮jl� ��Cr3�`0 |M�����p^�0�}�pe�}5�? �ta&@�g=%_r������
�^���.����C�	��M��~��{���.5�i���ف,s�K�5u��Yj>}�_ ��3a�v�2��-&�1�2{dx!������qZ~{d�K�g	yc �#Gc8��W����hn�bQ	���c��}�K��"��W:^���G�m��K�73��2U���9Q2���~�Kf߰�Z;	CY�B�u��K��5���UxݠH>Vԝ��KX����L�~(T5��xF���wH0k�Q�ŌJ�Q�,�k3��י�,��}I��Q�a����JL��X+�W�q�UKWS�BL���ߙ�
�������a�	�]J��yэ��y��DD���mn����e5\���_��1&|�E/	{����ѝ6ɐ�o�wHQ�.����;�[ �c�k�ߖ';���*!�� �J�YYW�߶\�8B�����(���7���ַ�=�ըޡ;	"k:n㳲s��_]8�?I��ngptP�}P�F˛�*Љ�m����8U7'��'�B�|&W+�'tpP[�*z�%QJ�B?�9D��M�`8���� �?{*ϓ�[�w^t�������q���O�j)�lIB�>���S�t��9R]X�[�%;�ῢ�;��PhC����JL�w��4��W����R���%=����P����\G�`�$�$w�M�~D��<�M���'�E˵Ԡ�t^��b��=Ά�Gɉ1r���^���{t[6 ��tr��?�&o�ὖ����'�(%�6�n?p�\[���/M��u�A���Гx(���	�ɔe�洮?��b�Cݑ��ۃ7�2c��l"ß"�~<�EpF>	P�uZL��0�:e�Hq�T��3:��t9�Jj���K	��}���iW)��g(�H�ō��kz��A��	��o7,����O8�����"j�Ēl0H�=����T?}��u��i����|+;_3OS��q�Q�wp�cY�j�L
��H��\f��L=��i��^!���!�؇ܩ�j@��ߙ��ѣ�H�HL�D�����~�,j��+�̕�L�6*�	K��<�B�f���݀����UYe�fB�i0��w�H`���m��U��W��d|�2���}����x��<��KryƓ�B�m@� �NV!�-R���@hA;��5���0� �����՝_�`&|����������Z�7٦%F��b�Ն�����]�U͓�+�B������$�Iﳍ�ʳ�'2���MWCN?����%�����ZG��Ab�(�9�j#%H�~(�����'��z&�>qUz�}V���$�z�o��Rp}��X������:���F�$ӷ=O	 �����g�UW7D��	b�w�Qwޖkiw~��	�g1h}o[0Jn}6��eA���(�\K�m,>>�˲���0B>r\���K`���X�z���u۽�a�0�d��p��5�tq���Ė;�f�!����~���]��B7�$��Е�&���_0�"������?�r�k7"�mG.
�^�8�����y��
%(����B�=fh7���l���Ͻ�z����(F
F�[*q�O��*(Eo����~I����<�&i�؂d�3��:�-V=��+@��Ͼ<�>�� c���9�T��³���]&��M�@�"��	�pQ����ix��uĥ-���)���C��u�+E��^���Q�ڵ��B=_l���(�Wg���$S/��S< 5�#�ߖ���L$�G<��,�?hu�%m@$�?j>�!o�SA���@ ��[[葼w�Z�
��JL�ԛ���pk��?���ԃ&����_��\:uc���% ���#e��j�������y��q�H�U��ғI?�p��L'��{|)��	�EsT��V�ћ��}�	]s���K�u���n�b�&�X6j���k1����w}7����}��Cd՞|/���5�A����6&���mL�\WvvkXN6 ��h�
@#���N��1���W�f�Z�~���;KvՀȊ$�^7k
L@�d�2/./��3˰&��\��5c�?n�4*g,c�|�ˇX˂�����A���4qPOS%�P.W��<�#Q#h�������נLF�:���w�u�K�y�/�
-O��� ��1����De��r9����r]��`� �	�(f�����Z<	L�aYǌ��`bB�����ެ��;���dtĴӨ�yv~
�w0CL�Đ{�zq��qa����z��7E;%!���u�nz��|5.
�|�gf�R0!Epk�,�C���|r�/&u�OE�)��މ W�(�;�W_��}�<�'x��Qdh�������l�s(j<��4=z���$����h��9���z�3}q^>�7^�mLr�4�QG�f�A��kNڵ"�p�Ԥ��Q�0�u��`�,�f����C7A�1���Bnڋ?^�?>y0|��a���k	�����ٽCCd.qr˵�f.I�z�1�o%���3+�^��!��M�˃�����fz�B���ȳ���ǿ��j�(~�zE��O���tp���(��Fm���K������p�?e I���\r-����>�7m�巀�{�|�x����UW�V[�^�VL]+�����b���M���{�14����c:�����R�1���j�u�ݜp��:�$#p\
'�������mr�=�X7^���#�	�>�h����m�B��cqKru��\���-ï��� ��+�aQ@����v�Y����<�m���6;)��-/]=�\0<�� '�(�#�RX,݀����`:^a_QQ�kJ��=/0��h^`�5Δ���F>�g�#m�/<M��-������ap�:v-a���o�x;�$���~��%<�����G՗r>�Ŝ>;�.N����	�3�c���3��P9�D<h:T`@h��*{�2�H�q'��MW�Y�)�t�%T��r���@ݱ�����hDh��-� 7Pāh$w��a0�I��Ӧ�fR�A[�qu������������E&��3W9�ʫ���T�X�4�e������n)@ \.����oG��K��c��I#Q��1AIɯ慪�)mV�m6����e&��%�	'�5��<��~�i=Z0����h�,�@�#�P�1��.Hg\E��ች����w�p�A���Qa��?LU���Q�f˙�K�֌@`��b?��._o�v�J_s=��3A@0��#�?��z��q�����\�az��{r���-+�F�/`�N?�&���}�ۙT0�
�T7Za��V(���R~���֩����u(��J���S�8N��_IN�����dj$���vg�qG4����ZLǤ�k����2�~�W)B������9�AeF�aG��.�8l��E9gɒ��L$I��b!��Ol̬�ph���F��^���S��Q��n��S����6�Hî8�b�)���7y*T�$d��7tA�@�K�u��-mv������5|�贋�'R �sw�s�/y混�ZP%W���5�n�Sȱ�������
��އ�|n�2�R`$�^�=4����%��-G튪��c
��3�3y�H��~h������'X��RY�j�oC��TG���ՐT������P����DY��)����ϟzb��~js"n�%.�\�'υ]���G(yN�{<ѝ���T���ޭ����ڒ֍����k�N�nq��:�&;�+����������*�=���(�ړ��-���9a���4r҄��͡��
�ջ ��Mwg���z[���t���M���D�y����7�'˫���%��Gۥ��d�c���ǤbT��g�a�/�p�������Z��%�p4Ù
eu���>}����m��v:���+���T���'��p�^
�vlPȋ����L�X=��T�A����ƨ�(�
�X(�U�9P�?�_���3k��_pl��-l ����$� �'�*�d�������â�7U�n{�v������@��i.�`�8Ԇ{!q��n�AP[t��"m@�Al�ȓ�����◯����Jѳ�e͚�担.S��j�@7#1�����I�3�찚�_���k���v��&=����@��7�tknȡtm�Q9�E�W%:�Ufbi���~�ͼxc��g�R�O�Go@�u-}��}��Q�vZ���p��r�ZH�a���e�R����Sd����~N =�h����g�K�̜͆���i�����t ����=?�gģȡ�h�҅�8������;���[�����dq��3�b���9�/��=���V_�����R�+�8S�ف$sн���!�}��!.��y���寉��'�@�/˳+s�7��dF�gԫ�����zR,{�Yf�M��5 E�G!�v�{c"|�kٖ�j���z�5�=GVG���=�ח�M�իWl.5��>��T�����Jͩ�i>��Fs�u]C�')����F%V��^!kܒ kt�';�����nܽ�������6�6��c�]ϙ|��/�gg��ȍ�a�B�du��WO�9ՍC'��wP���}�,�~x'�⁏N�_&;�L��
js��y�6��N��{��3�Y�hǆ���׬'��o=�ҏV�PV�fOXx�B[�����-<�N��U��'DGꍦr��Jju�k����9�����Y(���AmŸVyac�dk�Q�/]�a�R^���e���i��l���UR9K��W�j���b����m��h��URR�K���1ͽD%'O�>���`V�����2��H����!��r�DV7�&C5�sE'���������>�IqI6�!���Z�ť|m���D���Nm�Ծ�����F�!�5}�4g��òFQ�~g	�)���Z�����52�;��r��jmUK�b_糭f��;}��mY�Y�<e�V� ������4o/�_2��W��M�J�h;�f���¤�X�:{�@�}��7	ŕ :�� ��Nb���{a;B��Н@nl\.JGO^���no��we_�����;�&���J5 }���/՝��/���d�Q�.L�={�2���4`{$����=��Sn#ME#�i�g�ĳ��!y�o�l�+��@?�ڢO�I��$T��Q [�������qݯ�#��Ɏ���^Ǖx���Ky֡�7����\9>�e�ɟ-�~��(~��SrZ�ڸ..)�R���cEA?y��!o��Ӛ��/3��Bݯ�űPo:ύj�H 4���`}w���*�OU���Ǵs慣B3/e�X�k'�x�?)e������H�h�5$:�XC��K�����SP��3
o��B=��ط�Ə��3SX�q�EY5�[1���:~���'.wr�fz;�@�Z�dBS�_��WHMA@�C���oV'~���㪺�O��.����/^/��r]�?�P��L�[dF vH 2w�� e�A��9;.%� .?+�_6;��͆ui����χ�T'''|4Z��@�޼y3�
��wU��L��;���Ԟ�WBlq�Gu[��� �Vu��+i�7'(���5?��ń��OH���Xs��o������A��4���e��a�L�?Ɍ���2&��ы��z���c烍����Q�y6�uPw����I�_-Xd��4����%5j��pT�e1P^���,c�s��ݘ�dq�� c�*��B��ҳNl��~��R�� 	O@Y��rӖ�j��X�y���;>�4MF�#*���W�2�-������>����/��t�1�$��?���D�w����a��'��}�=�w�  ��B���F��I��p)<z�DaΨ�`�L����;��S�
?'����~���� ��B�������8u� e��G'?�c�ߜ`9����£/R9�}v�;t1O�q�=��8R��]k�%/���ybr��ւ����
��>��Lh��9ᡟO׿\;�џ���ۻ�];w<����ZʐsMf�M)�6����~=���n�]�ѩ��/�9���~�*cs�M�.R��J�jN-�*\<�<������&rj��||kj���V���5�"3\~��,+ �{�w���O�{�QZ$Hg��ڲ��G�.xN�[�m�&ٙ�	���z��L�+!)���Wr�l[�֦�0X��GyP���Q��
�v��6:>���@��J$��i��7z�h�Lzxt�m!����#�����SA��2<� 2�Nh�4GT�7j^ɏ�>c�E� ��!�~�Ǻ���f�S��Õ�cu��g>���4{��)��� 媫�Rr����P��R��ʯ~"%!?�{�8E	���KSO�"<����ql���J%3j~sT��i�MA��z|��`�j&3s9vsE�(n��޸{a����[�𓒑�>N0қ�il������Z���z=P~����o��F���s����,)%�sˮ`6���۪\R"�7^��x�?��{*�����������4�)c���9�xùE��x���t�c�y�wm��=W� H�I��X?�#�*�KX����n���	���d�ʿ/�RB&&����ο^z�;  �6>,-�x��j2Q��:U�z�2c�<�B��xǇB0�q��¸�.�q��6�z)[mgP����ǫU�&���v�1�ҟ�Y�!��q�C�0���g�Mut��^H�&ʱ͹OSn�>'j1r� 
8��c;��P��zz�n@\�tx��L�5����wR�D)�yV7Χ�����AZ�ZB�¤�hT�ǀݠ���ҙ�>�d�[�.-�1J��F�z6%�S5��:<�o��5��QC~�U���?V��w>YL����|̊�M4Ǽ��uUC����%�N���|��P��z������_OGT�	��:���8�H��y	�@#Et����V��ꯤJ�iw���/_���;�#�9�C�!S�7BD�F��\km�I_0
ٹ,�Aru��p��T���[���u�B̙�2��ʋ�N�d���s����E��m�C�n�i��u�kT𣝹eұ���-��e)x�e��
�cL��&��fY�3�	<:��� @��$��F q�:��h�S�RWȗk�ϳ��j5.*$�>�o�Υ	CDU��zj���;H�a���.�W�f�@t?�؈�M]4��1,W0��^>"��%Y?i�(.�m��}-&6d�q������ћ~N58 )X^^u뎣�edh2��%����+��j;Br���� 9p��4�0^��ġ�)��Z��3>�z?�h�����Y#=��
Y�`�<&-��CG/�=��V��TV�ח�$lPkf�O���B�)DvI��I�`{�5
ݎ���/L����mm�����͉BM1����J�:J��$k�{��h1��,��	G`��+�a��/�4#n��VX���^ F�cS���m�N����n����)00wHA�֠>4���s+��O�C$�z�Qydpph����;�}�"1����d���d666�n��=�Φj�{�:桴�Ow��}���o<3�&�pjH<��6���HO�uƬ ���=%KUѭ��z��g�$�04���'�LR7���u*M>��DX\6]?�"7f7����܀�|�4w�D�e\T��>LwHw��� ))%!�tIpK���
���!��t���PC7<�����3/|�̎��u]k�u�!�m��<S�z�]A�-�#)�/L��s�2oH�P=�R+�o�6w�r[�~K��l�����B�%��-� ���L-͖���å��n����S�ܲ�Z��ÁU8�|�ӲO�%e��+��&҄u�;3�{��t|��1:�w#�Ρ��N�f�od��*h]��>�����.h�2���*��5o~�@�Z�%ޔw�%؈��`�8�k��
�q}�[��/�$���J-�B��Gr�0��]6���yoMVV�w�_� 1�m�_y�vQ�~��M&3�n%�XX~_0N�:��?{���q��6� .�=L��*��0a���c��k�{)d6w��Z�d��9�\YI�1'K���Ŗ��`_O�$���u�ę�*=l����@� 0�*r-3TUt��G{�pz1t��1QtR����c{�V6�d��*�x*��\]]}����V�����h��.�]|�ҙ��0�yM�~��e�����{��Ϡ���_i�,��
3)l�����(oun��-���L����d^�F!F��;U��
�6�;ZLe07�ǥ��.��aN��~�Hh��	����ŕ��~6궟����ӧ ��R����$uґ�ׯ_P�V�?*�����m�rͰC�~�b��M�d�:&[ܔ���$���:w�y ������n��+�T] Q�!��'܃������Άw:��gd(���!�a�.9& �?��TL���I޳���]��֙�"��!7���MϽ �&5	���=JӾel�������y\��:2ϙ?�s��w�>3XK�ű~%����`:����A�`�]�+I-���'hk=�BI�o���k�a�0@@���������l�P���}�g��Dցm��n:I��Øӵ�HRU��C��q�Q!^^�%os�<K��É$jݝ?�����i���~�X�wJJ%H'����x,��)ά�-����Ϛ`f2֨��������Jh8Q
�g��D# ��ۧ��jlZÌ2a&C�ʹjt"����b��LV�BB�rv�p��d 0`.�}H;:�V��3�x��$���,��$4�'���$i�?�i��q�O�Q�	���-�C~dU#���h�;�����z�:��6��W2습���I�n�Y7Ҽ�Њ*�@�Y�GY<���9�5�>>��\�B��Ea��ai�Z��;��_��i�X�BFmcl4.js=�����5�ɧ5rO��	�Q���iHevq��(��h��.֢䈊�+�#�:I�b^�#�#��*k�6�/�Ě
��&w ���E�� N�q�l����/��*�E���jw~!�ԥ(��Q���!{V��NDP��9��Q�D%%s�c��-a�L� i�{��a�����K&�Dվ#u��߰����^�2�S����K�� �%E��]�����#�g���߼���k����D��s�?8�ϭB@��d��v3��T�WiG�|���o����E%��*Xrw��.+㜙�y���ǋ���Ә��W�*+9>��X��:�����{g�8T�AIBR��\�V���jD��a����e����N./��aה:]B��_ꘘ��@�����o�ѹ
�����'�R�����	���9֕�io)�.�E/��G�M���%A�xP������ΛJ�S �ﺧu2[�7����|��j��$E���`V�`����^���=F�����p7b_���<���Q��y<�"$�Ǜ�j����*kE���^�,/B{05�ʴ���z_񣒮~�8r�/�� ��t�$0�b��Z���j���=�|���{��o����/)](;BￓP����bH7������qUWlz��!�!��{{}CÁm�{��v��۷����_��"�W�H���l��ϻp,�l�B�OA�p*t�F��k��g�#q���)`���GM�eh�M���>����b ��y^���m^̇~���� l���1�}
t�!�5!��������=�q�~��t	`{o"��u�0����O��E��=�p�sW�|D��}	��}���i��w�
8҉F�10t�f�g�nz����m��Z
���V݅���D0����d̀@	^W�Q阰q!����Ie��E�}���
�r�^��EO�ma'��P�ֶލL��(�t,,��R����>C{[�r=}{Ĕ�<�h��2���A������`��8���t!�xd�5L���S�ݧ1:v��y�0�������|�����Eug��(��s��*u�՜�	��`������ޘ('����i$��0I<z�i����@��8n�OY���&n�+���u��&��ٮ:䥫��!r �&���9C��
 �}��xe�G���S��.�w8��J�p^\�R�o=G�_-xJHR�,	%�7��V�aX6}|��q��hU�j2l~^���^��5|���~0�,�}���|ŕ�x�r:B4�0��7FH��Z��g`�^����L�׆;
��(pYQ�����mJ��M4ݔt�X~ˍR���S1�힙�,�3&wu��[��!	x{9��C��Q]���*�;���~G��?�`�`k�G�0��e �u��s��0 �$lɣ��8�<#ﳙ�����9�e�4��R87_$��O��"��],'@�,�� ��~ѵ�iC#>JEeeL�[m�GNC��:�}�S[�m�� �..g�lN��\/)m8iἢ��r�(�g%\�����0.Y��좸��S�T![��F���% _�Wd#�cIQ탴)>XZ��F��~���� ���F)�V�lS�ڦX�q'��х)��Ы(����dIm �a4�G)���󸙢�(=o#����g+���P4���^�z�����TЋ�/���}�f.ff�\�v[��������i�[*[R)x�寋[�9ap��ȥ��^)�T2��4b��G��Qbf����pz�T�o�?6�_�#�#{��j���̻>R'ޫH�0.|i�TD\��O�����/����_�w���C%U�}�{�{�g�WF���B�p%8{�ڡp/ߥ��}�ϪTfN����ʉ�x�j�&PgU1/���B�b1nB�9kr��e����9)��LLb�
w"���C^���ޗsƜ{[���=Q��.ﶋ`^����T���z錡�0�}r/��2m�o~���@��
V���vZj'�{4�&���n�3�#�ָ鉪$�[]�n�]+��H����	,g[���EBMW�d@E\�x���LY��K��`���7Z	t�I���y�j�8��(^￧4��q�W�{�J��#�> �IBȽ���_�o0�����%� �}����/(�W>+7Kϝ�-���K����K�%�<�έ�2����ϱr�]��	�Ό��}�����ȼ%@@Y�R<::�h~A�}�m��A�)D,�C��b�o��Q2���������L��r0b5��d'YG=��,�r�}��[�u~������A�Sv ���o��"��qIK֔��ޢ
�:1.|<�[���ϡk�I��]����+����<ou���	4����C���H��L��x��V^�˪s�?�oy��%%0��4�"1�B ��eP.��6�"�U��T-Uҫ����G1�ˎL���;����k=�h*��/�>�/ @��B�B��&�i��u���=@�m���؄��8��A�����,e&%#��������s��}�ŭ����KC��<���[V�iO��յ�����}���~����W(E�k�~�0 �*�R�z�?��P�(q�����?;j�3�T�4�0�b���x��,Rl�m�V(|@O���,�x����0"I'=��&@�.}��t�'f(���jP��65�5�I�xo�\	#�=wP�U�D��R��ס_�~�}�?S�%�M����e�hߏ��]9Q%�������+�l�dq%U#��6�p��u~	I����i�20A����ީf%�$�o�f�p���r�V��+"��Lڛ
8�F��Qn���2{�H�l���b�y�4-�:�r�J�� X�3�^��0;���͉�������ۧ}x8����Q���m:��h��>(kg��R�׼P�}|
�p'��f�1/\4�&&mE?�_�k&�>s��h�Ʈ�J�z�	�0�a��7ﲒ,���{��������ӛ�$�C�[�j��ދ/!4��'D����v��<��g1�>�;�X���a?ER��L|�,�3�R�aU*YSØ�����"��bVg�lR������[E*���LUe�10���_ޤ����e8pi������p��0[�����߱I7��Т>�S3G/����'b/ڒ}������6�],��_d�B0��b�A�b��'9��}:�",��[@X������!>�J���/*"VZ��D�����~��ƭ̒���j$���s���Gr!R�LX�W�e��Ά�	}�c���h���U��|�R�N̠�gA	z���.ض���E�N�Л_EL��h�I��2�;¢O�(q���������1	�q�vt�|^��e�%X������O7N>^
����/~�ymg�.���m��uǅ�-�L��:��&����(�"�ƶ����
�OeeX������`5ν䗊 �X��~V��+rǆ�(}��`f����5��Z�
6�1 �d�Mb������hu�?��;	�+�}�"��RL$�EHm�6Lm���>����'�9 Ë�4����tӣ}P���sx�a&���\s_���8�L��z�}6����ս\X ��(���A�����>��r_��È)Ѫ˵TS���H�@��[#D��������)��g��H����9��;��_?z���恸w���It������+b��6u��H?��� ��uCt1�������V�+L�l��n��=��LQf�U@7cTTԮhߩ��ㆷ��ިy�vʉ��F9ߙ�-EU�u�Z��eX��UO �8У� �^��S�*�ף�s�f��6o��y�L{qM�(^}���mdܧ�����c���@ 3V��rF`b


�Ќ�Ru��FʁB�4ܻ[��*�sDFBdO�xp�������/�n�S |��S��@�T�L�"���D���u��Z�ߪ�U�3e��~���E����H� ��}�4�'4-J�����hak+e��!͟8� S�ު귤��Y�a��'�����ޯɹV>����VlӍ�f�Obb���͞w��Ҝ��C�s���t��'�!�O����V����"��bٳ�`0�ȔI޽{�����Gr�N�7m���0%I�Fj쉽�Y�;��e�U`MG���p�H��������si�?��9*,al����"� �f*�������a�&��O$�u�` i��hd9>H�����Y-4�����\��6M��C�����'�-ˮ�cW�9B�O�n�D����Bf>�%{l.�3/;I��,;��/ckf��פ ��a��3U�W�4G&&b���dhW�=���7�2�ҥ��ec��Si��������>�`�t��f�;����!)�#`���HE���"�07��N7�A=E�Q�+���a�D୰��8[�Y �s���ڀ�Ѩ�z�N��u먀�UO/�O��RKars��!���5x�Zpc�����$Xg)wߪ�;���R4X�� ��W9O�o��+�!kF���b��Z�o��"Y�ݼ��>�ǜ'c�o�u�:�����gg�bk�����P��0��uS������o��k�t��f -�Y}����_[�;�ٞ�dI�q8N,*@w*aS"c���t��W������8q�	�d1�Ҍ1��8�`ݡ[���ڛ0�i6���BJ
�8~���?� A�ʲ�%���m!���%&���
�nF!w��X�����N3���?}�N���=���8.�/�SU�U����w/�Eoz���V�e�=:W��Ǝ���e��~�g�%��(��(݁:O��80����P��LfpU��Mp�S�[��ci)��W�n��Ϟ_�\����ך���DE�</�!hau�,,s���R��D�e	zC�Q:��t!��d��&�~�d��{(���Z�
��0H��KcɄj��(�c�Ĭ}Ji^�(��dP�G��w?�80����b�o��}��%�@CUM��\G7���'�.��b�,���Bw���=�e�XRCT�.���o�����z%�4�i�-@(��K�~���;��E����̻wy&��$���+�\e�K��3�V��>WD�l�U�2xx�!�K�-L����PUv�u�Z.��9��с��/��X����.On�K����g�$���D�����zz˼] 	r��6��s�i��H+�:(�j��C2wdtt�<Ņ��G�;;,�G�rA��2Ɛ���s%�&FmsQ��ym�����a��
c��͏HH&�����k��9ݝ�~��z���.�ƽ�N����oNP߼VP����v��4P#`��Q�w؀V~��ZYU�	>X<���D|W����Tqyq��$�iS��k�)'��	�{�-R�H�]+!��8Tkݿ~�g��\�f���<h{�5�Xqxv��[u�w����� j,�GQ��K�'�("&�<5�.��Ҭ�.\��	����%��,z�" 1?��,�������)�3_�'z1�Φm��_3Z$r�\��z��Ub��g�4E�� ��^�NII)��$)���]\Hb�D>����P*�}�Ւ�()��W�,t����������O�(��F�� �j1�º�FFElX���A�(�F�#��\+����`���b�q�VPG���E�s�#���=@��M�����g��ǲ��nR���v�q�~��=<!z��r���q��9 "g`�_iuj��~bu�˳�O���a[��V��\wm�$���
� >~q��hO|N�cc�p�'��-&���h�YF����1Q*�3�q��M�77 :���h��;��6Uذ�Vr:�&��PT�@�4lf~ۿ���:��){l��o j������xK�ۏ�v�C��ی�&���п��F����D��)P��h7B�72⪔iD�B��8�����[ �4�ЀH���n��O���座?�;t\x���K�\��q,YZ���b.��E�q	���� ���/���f�یwo�'�f�k,�j=�[L<^��9��L�b��t(}��}G��*wϭ�gF�]���O$1�T`_=Hh����b� �㮏�'N���Ϙ\��c�t(�R_�����r���43N_K9�gŌ��72���&&�(��s�?y �5!�q��rr��^���q� d��E�D�K�j�x�꽵�d�A�O΂�6��nz0��1aE|�3��H��1�������Bکok����י�-j�Y�M��qh�y��wi�A�l��3Ѻ�@V�,�Ͱ%r�J�kW�8e͇[S��;��O^�|8�����"�CK�pv�td|<z���V�{ґPP���u�<Ғ]�+qx�k�D�0����\(Z�Ĝ.9 �}�׹�d�WqՆ�@yj�d����C?��Q�x�>ؾ19 ������}���Q$gPI2��^�1�!���s}��f��,$/��"�I훣G�;�U,��dvr.za�Q�|3U�1y�Ty����R:���p����O*��vzꓥۋQ/jO@�*a�p8�_O�"C�'4`�N7��9�{䋪���V4�X��O��,R��`f�)��¡ӳ�Dh(�(�g^?�W�r�@��{?��r��)Q���D!��W�>'��=+��r�I��.�.C��r���>�G�^�Q&u�j���V�'OFFF�Ws�ŏP`�OOOqb�f�ɭ�}����_m�c��E����z�еo��﷮��~�K)>�6�iS�[����\�=�� �ê�vb�D���Z�+�vP�c���כ�d�q ���ٲE)�����^0�=�>���h�Hk�T';���&�y�� ��h�\ -�A
v�j�]����T� �W�����B�cp^���	���x��@�CyY�������4v@��w&0����{zc�~|g�GVo,3��XBݨf�C���n�;��A\|���F�0�<z@M����)b��~�Fz��q�f0��0b}���k#5y��X�E���'�\Y���sT��h)���B�X��j�N�᷊�����x��}
�wО���^ͻ�"�??�TRNz�����l�ׇ�#�q�F������U��a���`#	p���A�����)���|Y 5����, v44�X�Mw��8ҍ�}�}���Ĭ�������6��������:^��������_�$��֖�yԵA2�&�Lo9�L�Y%B��r[���F�|y3�8jo"����~�WV��^P�,,V���T����N�(-FĐ]�t�A��E6�`s��[�.B�+�DSH"~'�	X�t�n����Z���Q|x�P�1`�V��u��Ť|�EX�lqq����|���#�<`���*RC�.�X<�P�#���K�4ىFw"���[�����WNU2��K���w�x��?;�?�^�j�4F����s[9��b��mL��H���s�������X���c.��[��"1�{ν���g3o�:�:6&E�Cb7������2Co�m^8�����Yl�{~�����KgAش����*�����v5 ��d�!aX3s8R��=ȕ�D������r��m�ڨ��M��r7�S� ��Yaz�;i�W�kԵ�!lk����&4w�6Wu�[�+[��F�Ƣ�Rs�x 9l�1����}�M�l�6�G����m�?0���󁈍���nʡu��,@F�K��<���Z�� c�jk�_Ce��4!#����r^��;o!d���.G�'ΒJ#��E���ӧO���  N{��?����)�r�[�}^0q��AE���┽��-s�Qu�L�o��AoG��I���{�PӢ��K{��7�J�P�W����G�T�q6a�un�Z�@�Y]��X��&�M�-K�5�x��1��l_a��#��g����u�(��/���<��8�����3�5� *�����Q��`xu�8f�m�����z;�5����ܙO��m�%�-�v�������LX#B^DD��r�>�̍W_6Z#4H�z��/��H�'�\����W�{-��؜ͩ��80���i���=9�N3p�����Z�$IY<���WPX�7j���$��\zL$��-�����Aj
0�c�X%��B��>�Ψj�np���E���@�q!���ѳ�q��K�GzF�]���}@�t�TO�|����wb�^jx%�{'��WbV&���i����o��hk�'�OBo.)/��KT|���nnBB_�c86��9�d^�Ֆm5�D�5D����x�C��F������j���a �X��F܋ƥ�q�VVF��2���w����,n߷~V��؁��k���\���9��q��Z���@��z��ZQ��77C}x0K��z�T�F�ϗ�PW<f׻X��%5��7��~'�M�g��\g�K�@4A��-,����5�B�x�m�?[�(�[uhb������c@��J�t�`�(�����E�h8�c�X����-o�_���[$'g�s���	zt
�VVz<US2Z��KP�G�y�&�l^t����K�"�]uȻO����a@��/������(L���Rc:!��*\8�7�! i�z,��h9X���[4�l�3`�t�j��j�t$��:�8Y˂�D3��|�ѹ����"=�I�u��N��Ϳi~�G�������[�Tvq���SΚbsur���޵L�E����ScM����SԂq�A�	�>@*��b~�v�AUm��j�OP�w��[ R{𯨪�.h"��*�H*D>�s8n�������O� �|`W��\��ڎ#v�ة��;̖����]�oOB�k��3���>Ʈ��W�o��V�`����R]K^�6�ۊ��~��',�K�ǸI�2��
>x_/��E�ѥ�E������0�<4-��U�e����?��\��*�H8d��)�l&�8x��8�����"�q�7r�r�Xv�.��[�i׳ �v��w¶Ԗ�P� �1�t�2JF�M�@?���2v�:+�|��^w}���L���W7�DSr���J��5aGI��Vҏ����u<�L?a��é�iy�r�-��o*�)�ڳ��_~~��Dcc�3�������H��q���u>�c(m�Z��'�0� 2.�S<�s��^f���}ܩ^�=�o� -��CQ�ހ����(�NH�f������	W�;�bU�A�]ߪ.m5�SP`uu��i+�N\�1��;0Cn����Hp�� Ή}�Ƴ9�j_�����i�Y��c����^Q�jZ�uVs�����W�u1���J�����7�Q<��B��/׾�׫s���Q(D�W���:7���ҍ)�&x���0a�&�,�)��姱x�<�B���Zpz�9�1�������6���d~'{~�U7�=��Y?$��	�'VhC��;)>�f�bv���ˀ��� krf&R�=����dW�Z$��up��%6c����>�~p'yrO/z�-a0`�����q��ǌ���'_��skf�W���/������al�&2Re������Je��@�ʺ��!@�QJ!��M?�^l<#{o���{����4l�M8�vc��r�-�b��⊤e����
'DF�w�W'��	�h-����Q���ٱ�MXS�3[�I1�Q����T��MLL�Ӯc��eX����xpz�:���֡�?Ś�s�������^B�z�3/�KbYQ�K�%S\d�=���ǌ5�k^��]��+�{-��jR��l�:�'��(�btB���� 膱P�J�K���D�q�[�����|��;��x`�))߇	;B�J~�3�:ӭ�I��N��^/�bDQ ���H>ğ�E{$W����?չTҞ`�[���=���� ���]]r.� W޴/����98� ��/A��^x����q$EP�X��6γ�\��z�k]j��'�A���ҝ$/y��,�1őՅ�_�Y��K�=6��zha�rob�;H=�j�d�e�$����ez:�Z��;���Z��jO#�O̘��q���L�Wo�I�����y �/Nl.I
�"W�� @B�@�Ízj��d<���zc-�ϠfYU$.���jm�g����ʦ�4˭���9�	^�
�^���=���'�|�I���}l<7b�U��&�o���g��M=��<�u��s�G�Jn|z���Ez����<ر�Է�y_
�C�q�rso�Q�n����k�0��F#��'��
5�*���g����?~��-(Աw`S���1 ���[^J�3W%�c1!����|�K"��]+��W�34��{$�N�@��)���s|2'�O� �`:~2qw�Ta�ww��*��yV�����c��"��Y���Q���t��g��7
������Q�T�+۫5�o���e�n/�#+�*]��q6��8�|�4<��ETd��`�o���!��Ԯ{��J��))�&��H�G�'�����!bل>|P�Јx���q,�D��1ۢ�����u��~�V����	JL��Y �)� vi��j�����?�+O�C��y��ݰg��B�̥W_�v��\����B�[1��5��#�À4��Q�������x��������U5s���bp��e����ꘞ1�� x��α$��w�`v��A�8�,�&�7�7n���mW��Yd?Z�i�'�T&���-��������B+�������)؟�7D����p�*J?��������+��&/�Z��/����cM�C�$$�H�'=��+g��H=�S��^7���&p�P
?�>^�[����Wz�:g.��jk���`B{�$k��s�`�ƽ�f}_���^±�OfO�m�����,�	�`VHh0�E�%�e�AR`��V._F8�-#q��|�7��v(G\��T�cd��DM�ɘ`���J��ggP�22�s��y8�@�L��>���!���3뫧00��ǅh�$�GV||�)�>��m��U�^v���N�(�~�&���N?��׸�	#Q���R������Id���>z��^h�A��{@ez9�ч�2�h0����赠�b��Y�����4�x /�e��	���֝{��%�7!H��X�Jx����~'������"��L�M�ZF�m�������M��|6NM���N��^ƍ�/�c�kQ'�r�WWMnE$��c�|\-�d������m�����s�G7��W'h׌!g���u��Jd�ƞ�.�����W�oK�	���^��"���6/�(f�?����g�(O�+����pKi�&�x�^�&H���CI
1#,��]���.��H�;�ȕ�If�'� ����~�m�J��v�h����ѡ��(�G�t3�{�Og�I�
�Z��A���Nz�`��%ߊ���r�_�r���p=����w�;ʇ*��۷k^tI���~�[�����߬�#��?�T��v���%w�1�WWĬD{�F�c$1�����je�d�[�M�U25���&#�~�|g�Ķ�Ċ�B��U��g1��Z 0�*�c�'���>�x9�)}�&&}8�i�;}
Vy����T+ol�&�./�Z��33^[a�u�
����v��H�e�Q!ϊ7%�6��(2�׋�?�zpI�Xh��{���k�(I�G���,�>��_ĽO2<#�w�6�8�'���AW�7�dy�W�9{3���j�?�|��C�����j��R;��)� ����$:V��\�_C�-�T��Q=��͑��V��v��uE?���7�=�5F+�+ȗ2�'���iSTm���zN�,��$�A���Z�I0r����V7q��˽��D��{k�)��&Z(f���\`!-#V���\�;ρФNĖ�J�V�/24b��bD�k/�3��F���~��@-����%��~U��jwO~��9�n�۲/X�#F�AŻɂ�O�(����ֱp�~7�Ć���V�!C���;z)�t��R������*�OLMO?���n� (�"�<ƺ�}75*��Dw�M�1M�З!��x���Q�:۱�J��[����:#��(83Q�����Qg�4k��+�:��iL���h���x

$4#�5���.��j\�{H !��C���dS�)��$�v�G��݇z������a�v�v�O�vx	�O�qQZPc� @�P��<X_F>F$�vm<�>��6E3��.I9+��n�:��b��|~��4��{���dl��_��+H��Y�ݽ$��j5������_.��C�r�Cş3m�g?�/��3�@��9�X}��<}�׍��=$4HnE"���}z�}�e@�fEw�T��ɡ��P��/�R�XC}Z7���#EO���#q��K�Ě2�+�`\��֜��>��Ч�� �'M>f����D9��e��j��<�s���k��d9��0`��d��mEkC�P������b�3fXY��Ć!o=~H���(�'Ԓu��]�55�9�ZJ���p�
�f<����`}h�W
�y��s��D���#�V��<�
��rd3bp�8���� !i�D��5�^�	J��=�@�9TǳAu�R�G�b���~����7����g'�'zn��c�1�"�L�A��@�x�WcOlUc����}47���5E!�[w��K
����ء�M�Um�z=�C���cP��Q�Id�8��S ��C{��I��5�R *f�}aM�wK���������i���Yt��*"J��)ԩ8-Z��{QfXc��U��g��,�s{�<2�	դ��g��������>���/(v�e���<x�?���01�9��V�5-߳}m�R���+oR=�Bq��ԨsVO��W59ɀ�i�G�U/�$* ����h�}KѵC��շ��쩸�~&&=+줊U+Q(7.��(��s%�<�p�X��`�f�t���~�� �
?v�hKj�_<ZdoM�\� 0D�NP_t*���o~������h�}�N����u�2��	���[{B��s⭷�)�]��Ϸ;��c��$Z�V��Ld �A��BoTt�=��o�E7o��Ђ�ܫwv���kn���,���Z9�Q�^!ׯ_��c�h��+��@ƨ�B��i���������d��T��� �r](<(J�A�c�,�^���Z��.���� �Φ,U��T� ���5\�����g/���Z:����}��?C@5�~]��Y�����n�t���KV<��eAO>;����G�c���Mh��Y�P}�*�W^M�O���^�V��VN>���~"Q�m����6��~Ÿ�t�ܚ<1��#���d��'�p,��@|�#������!fQ'7�9�i-�C�\%�Ê|����������@���Q!�9�S�|"S��h�W��A8���P-&,'��0ǎ�:�eB���OT��(�����	�z*9�=B|Ntc�
��j��Rg8)�lZF��e��ܗU2�(��n�v<���Q>Q̖��>�.̥���I>*��lE�3JΕ�n�^F��>e�
eN3?<]�u�';0�li9E\]���Jl��,o?S�J�}k@���h�M��׊���<f~nn�w�|��~����D����j�E�02��k&u{G�GE)_������HGF6.�Ы����%Ŝa��daJ��Cr{j�/��fM�d&�����q}1˦���Ɵ��KZ�P����zB�I=���n�n��Ew�{-���زYX��'bK2�"�:�rh���[���ѿX�.}!_>  �$s��J��~^��m��-�^��Ǘ
��]�VY�DN�CL'�B�(���F��m���f�Q�,C1�w&ʠ����n>�������,!��|!TTZ�o�i�J:�w�B��6�&�u�Һ{u��ӽć9;ur�-=N����[�l���^��-Sd���߻C�� $Rt����M���Ԓ�g�?b�:p9�Z����x�%��?M+}+/�m�l���@ByT�1���ܨ�1�]2�((˼xV@קB��Z��.M����Ć��'Y�4=�;���-0�DN�����)`����s�Y}J�[�"�J�����ߦ��ٷBi�Ge���4J4>qRM J�������S�
����v����t)Ӗ0�W�g����xf~�\8�]&���c5���q�������E��9P´�(W��_e�i��ݧ��P�v���׋�c��P�2oQ�y��[F'7�џ���}�{w<�B[�oV(t��w_� }�c�x?�dI@f�E���-����d��ڏ�����n�#��($ʱ�m�b�/͎Q3_�%�� w1�x�NJ�A�'gg�����I66D����ř���b��gk��l���z=��o�����ӕ ���%m$c��z��~v���Y�Y�h<q[�F�-b��P��ƋQS���,��,X1��۹.�;��Y�Hmb���� ����6*`w`�)�q;D>�*�dWY�[�h�JP�'�)=�e���J�]���:��Fۺ�m!�����9r�4�υOE���|ۻ�[�~�����/`�Y(<������.&��ӻ�4�(��)�tL�B�v���3G�x*�ʮ@ā��#*����e�h���Xѵ���W��p�ʔc��y���N��?R�_�h:���W�^�����&��tЃ;�|��d��[�>�Wv�K�B�=!�б�+��ޖB�Dtc��d�~1vڔ4����q�\ɄZ!�P��P��C�C���vE܌����[�>��?�R�=u+�F���b��E<�i޷cyq���K�G��`EZ��Y�#�{'Bs=���)ؔ�H�ϚG�v����~U����ֿc)��8���#Aľ �ZD挵в,�>�-ጳ(��S\b���������c�;�8�s��O�>[7���	f��]�(-�;�4⥠��TV��
躃���V�кT���*�<�%!�rJ��kb��EZ4����8���L�y���>�?Q�;.���_��K������;k�~�t��q�����C�&t<�2��<^V{�w0��{s{n�u/�a1߫1/ #��?!H<��x�aL��%p��n����#n�~��64pB�Ğ��T%�� ?��H����Zq)��aPW&��ɭ���6͐�� ��]Ő*O��w����ߩs��J~q'pw!G����X�l���T���l�2v������CH�9��|�م<�h���'��c��*۫��~PnЩ8�\���u�Uvȯ��}l��溠;��j��Y��JLG���ø����T»�o��#lq��O����9�Q��v�<V�7�L���9��P��੠z�Uu���sʈ?v}�|H*��Q��lm$P��nO}�I��sEr�=tm<�(�97��~���>^�~b.[L�h~fkk��w�
�@4�62%��t;Zϡ��z3�S�Y~���&�*���-���ݐ�B/[�"`�?���3?��ayD��~��x��۵��j�X�Uĭ@>d�/�N��:Z�ˣ�̫�V�yR�K����!�+Mվ�)>>��G7*C���T@�$���񐸫��wI� R��n�͌�����rf�ga>ɠ�
�B�Y�f�7K��
G�n��\<A��Flx�Ť�nA�F�bڙ8��]�������!�'�q����}��U`S�Wx��آ�9X&-���<f1��րQO	>\'�����rbs
9�G�y�r/D�z���G�*���xĉ#ӌz4B)bv��l��}'�=<z���#��-�r[/>�m`�4��G�eQ��V�^��������)����S`��2,b����w,, �8h�;��r1靥ooݚ�J'�3A�My�fl���C�)T�Yq�ù�P�ڠ�8x���x}�]c훪�l�1��T�['��ߕ�z1��z&�<33D+��׷��2Z��`Te!�y��?�*:�����5d�4�6���I�Ige�ᐬ�܁,��(��c�,�����O�Hw�R�]��tw7Hww#R� �����"9�������#�������w����y�9�N��r18�e:�&�pZ���g�6�+B�ǟ�܄��:�+���^�޾�@K��+t��1U3lv`��D1��|����v"I��������W:}���QQL`�V�����H	\�WL��Q�%!Bs14�����n�_1:PD ����Ë'9��N�!��-<������/U�Ô�S�YBt�U÷9�JV�ɰ�$e��e���e���$��l�HGs5"��а�{��,�C�70��BaأL38t9(नm�e����__���o��&�� �~5�$g���'S�!Ǥh��1�����2S���� �i��ϔn���zO'��E���a�:�F�?^�B���Qn������XJ�T%�`�¢��C�!)B�L��J���RDEXkվ���3�0���lْ�w�3a��x�����y>���9*��E[�n0��0Is�!��̔���t*�����2B��0<*�P5BL�S�r5l�{��]kcu-Z]ƾX����O9���Y%��,�t�!��C���vߵ�h5+�*=�C��V@�I46�  �0c�$n�񶃥&	�,�$nT+�0ڶ0���s:+�� ��A��y#��?�@zrP�f�m_�۱����6��5vk�{n�?�Nu��|;���" ��(��X�a\��/xRZc8��d#�A��Kl�;p�(#%�Z2��|����鰐7�x����*v?���@�� �2�Z���q��Q�/�`�Jo�حX�U:����-D�ʙ�P^;7"�7p�ˍ��h�g0�%��%$��S=��j�͒��Vv�k��o�����y2�wiku�H�zF�A���_1���D�~󇳇��G��xbT\�����'�	��3��!���Q픝F�<]�ri���d��5�;n�]�<�t	>(�/��?v+���}~���|u�2Ξr�?�ޘ#�-��	��gI������K��xQ(�P��
�8(�1�di�xCt�s�n�>��iX�
<%/8d+fd+��(��2��q2�:�U��܈������R�:C����hT������LA�'F1Q� %�w��S�Efc90�gfS����}ϟ0�I��\l��0����`qN��M��f�i�O�zh#֭J�6�8�G^[H�1�1DB��ɵ��ř{~`a�y�Lу-Z,���F�b����i����H#`6?�7?`�r�qH���T�<�\1���匾�Y$"u'���&�ǵ [4�0�����W�)�H�($�����	��_�[5��Q1~nz����@^���O�B�>87o������~��*�jug����H\�9�x®��Co|r�:����?A0�9�P��!��J0Vo�EBԩDб��D���L��!sܻz��Ǽ���v��!ߺ|s��R:N�;d�(`�,`�C�)g���+ju�L��!�L�5�22�0G��c�v���ʧ*M�mU����d���a:����� ^l���r��w¹]?!R�G"����~/Lvqh����*-�~R�EI��R�Z�)x��5�]����,�X�
Q���\.����L�G�H����{~O��N��öiRUJ�M�r�o���۲����A��0]�w�7����짎h$�]VV!/Q��篿&�U�Hz48��֍{���	WH����	)u|�^��L���3H��lk�d%��;�ʛ��]�����zG�l���S�}�itӹ2WUd�]���I��d5*��)�O��	�"�d6�0�#��m1;߶��%!��q���[@�4��%cf�Q�G�I����i:6�-in���V9���3�SC zZ���e�Iϙ j� +L��zH�5��G��X���EmӔա�s�-.�����:S����������� �iBJQ�x�
�����|NɈ��]�Y_�`yϣ�X���E\�j������,�#�}��vп�gI",�=I�c���`u�O�L��x=�q,��ʔ�����8(@�yb��g<[��ԣ���{-��~�p�͔uR�\��\�a�*�\�0��B��__!d�#o>���0��r��q�����D���k����&ѫ�S/
x�[��<��2;,�]�b�L'[P��4B�g�C{�?���6�G�3'5.݋x��"�)��b�{w��ٵi�@U��9�KJ�7V���+BM���I�Z$O��Ó�Lg�v��X|���"0� F�'O�n'��AX�����/�)�����`�E���b�e��;�	�N�S��q-F҉s1�}F%��'/�+u�A����[C�MЭ�BZ��Kz#N�qm@ǆ��F�����?�?��lwJ�`)�9�|c��>H}\�C�ȸ���r!��|?�Fp.�+�~���ǡ�sr��9:�В/&����CQ��|ۖ��A���ӡ�֛������!�o�(��`\>�K�hx�v��������m��c#�����T��'d������Qe�@<��Q,-?�NT��t��|��<eQ۱�����O(�ù��Խ��A,��A�d�ݒ0���>��\X��I�>q9����a��s-�]��>�ߜ��	 =���ه����7{TD �~ԯ�F�>�,
t��)��ί�2B�W�cóf��Ko�Mr�8�y�;��N7&`N��)eH.��c!8��~M�	�6S���2	��wU?���k��Rj�W
���k�����@U+F��hn^���� ������W?���VJ .�ґ�!>-G��g� ��7���->���9'3�#Z�����s������a1H�hl�z�^��L�^��d}��I�/�������^�l��ò��_�r�WP�g�M�εujn[�Z��J�����{m��\����d�7��*4!�o�iG%�3b�Շ?�F�qZ�c���*�$�rՐr�~0pq�ؐ�,�m�{��>q����5a/r�K��
Ӓ7��鐷���-<��uޛ:m�γ���J��;Wt{E2��|rU@:�,_��)"�YJ�>S���>E���&R����+�ۻa�(��S�+�\�}��߸���y�6����o��%`r�i��5�^�94���� �����k��^x㿶������S	���JB�~h~oTa����ߘ�rԀ|�����? �����7��Ch��Ͽ��ߜ����d�{��X��1��wē�����P������h�+��ZL�\$�Ն
V"쓰D7��X�����p�n���k�8t���F�:*�: ���b��j�Ԃ����5�b�\��_�y���׃�:H��]�}�F.dm(��߲=E�8U�{��pԐ���Ó�5eZ,o����k	 v6|3�(�$Kn?�PS'���s� Kx�
�m�`@&�%Wwq ��',Y7P�5�>t�`a�����$�ԅs�M�3"T�����˼�yToА�\6�$�e<q~�Re�6U�1ִ�M��s>@^n�Dr��Y�G䐓�  ֙����%�YJ�;�2��w��d$�=�Wu�-�U9�a�/*7�&��N�_�;�u�"-h����DCt��bc{7Sʫ{�4a��!~�3�����N��9�슎��o��E��g��Ц#�2^2f>�I���e�յ#A��c������䎿B^��D�Y�c#*S�*?���|��RVml �-�:��=���a�M�*M������F5������������5��������ߋj��r4�)����\Ⴟ&=�\�8R�l�b1���C�ox�ҽ�&���)aG�U�>��W�J�=�v@W���(+�.���CઆW1�i"����E݌C�Z;B&���/n
�� �-Q�NX.i����%¡����헰��� ��� Գ����n�P���zߣfn,P&�.feE���|z>�~��f�M��2��>�U��cĩb�������|!�>z��-�%wH�w��p7��F�ᝊ��Q��JFA�כ����N��y7cX
�K�0��pR���w��\oW��O��R�	r���i�ԏ�؛��k>���9�c���d�a�^E�s����B)n�8I�t-��:
ȟ���&u���r�-��*���
��;�)�Ƈii~��,�� �GqD7U���Xû�N�l��:�oc��	i%���K��s�W�(UKk�L ��MlDCp����*��cG7�����CN�G#.TA>���2�����/Ty[��;����K!�PU���y��P?��¾�ƥ�~����ss����E��9r����N�yd�0�}���t~n���c�?�*ȍ������_�.'�"<�=����\���F!/yZ�*���U{�*t,��vYsv�Fn9o�M��������Ãk��qQ6�I������7��M73=UM���{���Hu��A (�T�b�� � ������R�&�)��0_n��x7���za��d$��q�Ԟ(����;�����ǃoW��&�	A�ikvFT��8��K�����HE��a�cݥb�3���_3�a����.S}g_���"[<J��^X�d����M��	 ���N�������bu�1�?ɂ+Ⲿ �e
��.���*T�e����z�:�p2[�Prg>	��01�Mt�aa�8�UhwaqG�;wҠ�-}�R�r��� C��	D�{{ �u����G����D⫪M��aA��������A�<q4���Fx����y�s~s��ّIu$���{O�6�V���-4�X�tPu��gqM�{�Ԫ�m�!٩������4��-w���p}�E�;e�����L?\�[!�����۞�U��[>G�q�E�$��؈�?���;�0�����Hl0~Yگ�8\b�ٌǳ�v6D��sJ�7���D�q��=����qW@��.R�A��6�2<y�M��_��[W����x����M�9}�B��[)��9w����5 ��`n;���|b�박
!�To�S���`2���Ut!����3�� ��x)��k^�����N���b]>E��� �Я3{	08e����d5��B����Q�iZ��l���!��`�2$�x�*��+_��t�M�e�t>�QZT*�j:���r�Ʈ�~j�G�ģ+����1����$x���a��Ỷ�t�'^$a���r�A4��������):�Y��ý��D�͑��n ��g�U9Ķ4�C7���&���H��Y@�Lv��8��y��2������:���͍�N|[l��o�P��KQ�*��A�\ Y�9���Xy�D��{������܎0�O5��A�F߃�I�73��~�m̶W��03��g�N�7O��.2F9W��m<�X~|�)PG���4�18JFA�U�n�.C�~zc��q'��L����R���O����L?�����R���"���Z�����A� �������f�ޔ�r���� xGXAygs��|��~�|Y�Jp�0����c2����}�A�B1��y��<B/���������֞���dIo�J�� r��:�i]����>)gX~h��#��Љ@=@�;G.i}C"�,��3��[��?ϻ��Pܗ�]A����~�/5��WoG��<����`9+P��s1�	�܄I���д�ۢ��m��N���F�pt�?��I�#U.j ��'
q^@�?��ߜ�l�uS�ߪ�;�խ����$޾��h �{7b�]������lݷ��#�ly10H�k������2��O/�G�,H���To����k>QQJ9 ���ɽ;Oq�4�oBL��Fku��L�vgW�~�#�R`��K�ayoJ���&��j�Ow�K���h��6����m%�_y�5 ���{ǫ\ԃ�;��������ͫ��>��� :���J-��t��v4�`��Z�76�������jM� 0ʓO^�����g�[>{<�$�F�I�`?�(�_���Q�����Ȃ�#R��?����Su+/�BZ	v��M���=�/�r�ڂ��0�-�a��)��- ��߂���xpAN�]�����P8Ғnag�Eҝ��AAKA"�E������;��n�/���.�ŵ��D瓀6�|�L�I�"����(&����}�Yf?9m�v���O�)���8�ٜʰk,/�8 �t�xMH����N;)@4��dܵ��%�X7�6A����HFFi ,��V�k��`_F�oʁPE��셐d�OlLw���S?��1�3�~��O*�}n{|�� ��;-�P�d?{´~�W��S���O��&]?��0�:����a�}Gߴ�2���.x��ŷI{�x-�'〷g�/�51tB�&2}���N��+s�m���!R�u�4���R�X������I R-^��������L?����L �˯���I!�d��E!=6���@����rk�¸�2��u�QXT(/�׿�_ڰ�(��7�+�e��������G#��+Ĕ��[��\7oo�-�M�S�p���C	J�-�A�}҆GaT����D=��79�]?�,g�#���,�v�G+L�;f��u&��u��M밭���7� q�ٴ�Ү�ϭ���>�1.%����wd�6��`$�N��B�k�Z���K+A|�Kd]� /��Ϙ�X��O�9�����x��@5<�g��|���/{n�Mf���Ӱ�[�)�:x1�:Ǜ�%�c��p�'Y� 5������xwz5�jN!�Jk{�V\�a2�����%���MQM�24C���qMXR�wP+����`���Կ�c�SKl���R��ʜ"��R��q���ִnʀm�?����o�gc��͉'=��^5�$�h$�f�#��+"�������|���dj�y���<���r�g%���@q�_��>X��K�i�,e��i�웦��5(5QQ��ϯ������m�PΆ����Lt�,�	i�� �pg�����,
��YLvu��<��$�U2��1�K�:i8u�� ��cA�<x�T{xu�-��V�{g�
�7�L�J��x�ߎ������^���PW��]\�r��Z �w��fc�ނ���VE��;ʡ[p�&tb),�C��7C�v�f��C��U(���P�vqZk։A���yçc�C�Z�1���)�T��18�6�$�
Z^�z�f2h�'cP�8�!��~W j= ���c%��ni�6 ��D��ѳp4k-�1���Q���
'"�:^�J>I����LTċr�8��`b�bC6�o��8���5����#���;L����=�@��w�w�1���aҭ!Oj�|�=
������0�2�>�J� �,w=��t���Ipp�+����׫��bv5����#���Ի�b57�#�m�P8p�Q&��TGM�X �vɥ}O�f��?��d�z]N����9�ܷ"�HI+���%7�t��r&=�k��ߒ0�K�ӿ���'4�?ֹ��mL-,�ుi%Q���6a���3�u�)]�ݕ�U�L�")�u�y���IW����Q2b�/�"��Yfr�/vP��>�|����D�6��Tj�Q�lpL�o4��Q���ݜ�z��=[��e�c������Xu������� X���2׎�M2���V˓�R��ŉ�&�'� c�?3vVb��A^S�����EJ<i@e<�ő�β���cg�x2��7R!�W*~B���U?�����ZF�_Gx�4�y5�z�_������T>Y9��=���s�����(��u?'���A�/�F����!�S�H�����a��1��M���U��a�ٗVl!���ʋ|���φY�M���
ȇE�H��-NBĿ�+VC�P���g� �'�s�g.y����tM�~� "�Q�Ar<Hv'��E��p�n�*¡��w���⯮�R �?=��8и�&��gK���2��=R��|��K�KJ���_ŻVlS�_���!.����U�j05���q�� �����g�)��ۭ�˧r^=A����ro-��-*�m}�}���7̲�=A���P�S�W���e)�7�����^����ک�B}6�#��s��Wܷ����[�߼j�$Q�&iez|+���f�$,Y
X^7c ���D\��k��7e밀-��X�0�H��.�q
�������/k-'���{י����T��D������N/���X�Գ�����Tg�<8`⥄<r!GC��U��ؤE@��*O2\�{:x�������L���+KY �"!͒S�3V�K?s+ ��6<��ʀQ�Bݕ�2RZR3���{��AIpe�ş�r�L1�� ����-�~��Z�'+�M���|�社���/��kⶱĈ����\����Ƣ5p���uR���x+�� �Ҍr�r�'��v�n�t�l%Z���64��E�T1oDC�4������om]�Y���͒L��]��g�38NJk��J��̄"��]ȼT��|�\�s�������Ỵ/�4��$��
ʈ�X�aZ2v:�����Jfp�Qf�C�z����	���R�ƟU�KP�;WQ[�������� ���:ܭqh=�4U|��(�r�{����&�{���L�&��(uF���&C/D\y�6�U�� ���g�X+L���z���᭒��hVٵ��Ac0�p����x����1U�l.��֠�?K��@��39�0gn�W&s@6����6c����@�G'b�m,4{��`[��V��zO�R�]O���N+��K�<U!�)CP�h
iN�-�f�c�Km������j�}:�������HS&�z=UTX\��A�n��Vcdxqw�;�㨋i;��S����%���������	�*�K�M��P��ˀ��突��;��w�o%$���\@~�|\����DD��r�_ُ}f��6� `��i�*ve�P�H�U�2��t�*	�} ��^4[�f��X�q|�3��$�c`����f����o&dw�M���p�7��:��Է'��J{�W�ߧ�ܝٟ�A!�Sk�d�K�|����6�U]�_�w�W�#�f�a���Nrv_���@34�1�N�q��q�H���i�2n�T�;� ��_��'ǻ!�Z[5��.�짋_AG��uM]�'Ĺj;3˖M.n�������
��9iH�v7�8���S�k/�ݪ
3ȫ!\V�ɺ
�3���2W ��88�Y�
�q����y�$x�ĂFfg�=K���G������ޫQ{{��E�ᄎ��_,�͛NM*�[�P��
s^��V��'*Av�w>?�![���8���!�P1�v�$&�=|-��.�������J����k(5,m�:�A� d��@�f�j4iZ�ܽJ�p�73cc��|::�!؋߱Ws�E��ǋ�c���mһ����TΈ�2<$H�d��soW�0��	n H���!��7G����ƴ�8��>>��7������kXką^��U�!��Gw_X;O7��\Մ�j�J ����5��U�Ѳ?��oD�s!}^����^�_����$�L�^�����i%P��F� C�+��|\�ZJ$c&��n���9]H�V��A=DӸ�D
:����WBi)���+_"�u�&81c�#�l��CKumb����m58]
ǐAi_=��8�v �o4��T��f~��T��a�=NXVf���_��a���򚻖���QHb���fw�g���a��Q\��씝�Uj�2�l
b�>�Mv�u���f��o|�_����W��h
p��&�Y:.`�Ba�l�	����p�����l�` ~R@�x�i��,���Jg�Yr�ҕ�������#�p�	��؏�J�2����m0�,r�~"��oC�b�$�Oic�
{C2������Ex���6_ԉt:_�/��NA�jiο��D�2�������"�v�!�S16�C�ۯ�q�S���9�Rߍ �]��T��ء���r�os�9o��
��#@�Z�r\��>Z�K�@Oݬ��$��{9�V~Z�e�W~����N7����9��r��?#�s!:g��������L�Z!`gE4�x�)\� �V�Y�Ò�&���~�����.�1U�Yq����\@��en�ln/��%�/~���0M8�r�4FB7��xG+$F4i�=��yMM
�;f����z�@������ ��׭�4�H������Ͼ*��w�^���ى�@�!���W� �=�N�����J�m*����b/�������������n�t�PH�<d�wN�s�%!�F�=��P*�\�kU|���L�3�h�R�)���P`��:�#+>U����">Z";��\[Ge��ư;b8V�-/o��5��e���l��籫�9��� �yS:e\
I���PJ�G��­��C�3�V}a��b*a@�.�~�x�Q�k�m�1d�7%�P��ܕ��>�����,��� K鮛fnG���_(���B�_]W�>�S����ŏ����s��6]��OZ��5���z�Օ���,�����`<T��gl�Df�|j��$�W�.{3.�^	 �b��CT��E(-=�l\�(؅b_���	�^ޝJ�@����Kzh-�w�� d�����I3�����6`��lp,5߃�����g_&�6C�
1!��M�ض�^��`�`��O8���'ݮ�䊳f��-�.<F�^@u�[=W!�~���b�'^��:��b���{.�ϝ��o�w�o��>��eg�z�����Z�Ð�=�ݧK�o/�2��S����v��7��;��[U�V�#HT�a�O�~Ũ�-����$���R����Z>:Xv'r����n�)
�uA�^��/� �zl9xn���p��G17$=���~�y{z�f�G�Գ�ij0�kթ	K�}'�z�;\Z��.�쏰e�d!-Բ_憣���6֦������%���0��	��  ���f�螮�1��Gt h�&h�nx��ح�7}y�Ve-��ϼBTs(����Z�1)�
x���t�����{ғ�Áiux/bR88�F![8�#�*���������� |Ej�N���ܾ�Q�'EuP����(�a��z�b��.��@�|\w�a��9���{�吊�VS���������3B�����7�}�8��2#�P@/2�c	��u�ɭ+UVD X����˽��� p���>��܀<�^����`�]����)����ym�{�S�Bj%��&��en�åĿN��G�@���4���P<�}a�Ȏ�?�����<:����_�E�V�T��Pd|�y�����n�f��r�[D��@#�sH�ܗ]ǉn݊�,L|����ѪcLD�ڸP2*��!�jۡ�W'��z�S��w�Iq"O��I�<�(�C#bp��/h�dv"���MP����)���f۹%c��-��X�q�L��𺝫���$����?4��*��S���Ќ����g3�}?�_M�~�6(|�1L)�`�\٥w$Ү%u/�=	�x�(�@�������n~���
���qj�qWBZI��ѷ�zG����Z�6^P3/x%|E�r����f����������v�mЉ�,@�M/���Z�a���؆Ǻ�Xnn��-7yKul�]o��^�?���p����ܽ\�3��S�����gI�s�O:$��6\Ȓ��#��n*{�wfbL؋;e��]���v�s�\�Sk����.�?��R�Ĉ�5�͚�\�����ƙ�ar]� �yc}-:�C���o���J=�F���o���x�&��j���6�F�N�.��uR�#o1�,]��Y���r���4����`K˚�<��S��BM����zo�N�[E��.E6��X:�2�#�N��hg��!�G/@�����w�+��#�Y;x����ؚ��VU������!-�	�u&�Ƅ�`�j�F�N�ӷ�"�Y4���Kt�z3�q���q��?M?�����=U:�Uw_��ERA:��np�E�d����kK7Q�m��=���$�*��Z%|e+��߻o��`o*�1�g�(T.�V��m�����w��^7d���u�W��%����`���M|���k =�����;�����������Kz�����<R�E����N�|N�mjW��u�~UP��\'Χ�h^�1�5[��r�������;���bo���jxG}��u�֣f�6��Xn���a��'ܹ�3��/ex�����:���w{O�2ϛ��k����Ҵ��pL��� ��*��m�T��V�<Usb�3|�
/ճ�+��'P��<�A=A:�O�j�O�XP���?���di)�y�#�3TB%>�	~�u_�V��!�ʎ�M�h�@C8;S�LV�V�mA��Dr�KnQ�/�aZ��!]KD{v�&˖���t��`I&4.�W��@MLӸ^69,����G�n��2�~;O��4�yU=�TP��3���mD��/��h3YQ�53�Z�ɢ#6p�6���8kAC��	Q*�U�=����ю�*+#��nR�5ҡ?��K�QQ�`�N�����8���U�����@�^�Z\�k��\P_�O@\�e6O<>�{N���^���-[z�yVj�Gv�k�{����j��ǒ�]\�:�'�Bd�s��B��&��w:��o/��PSL��W���V�-�[�n��m8w��u���\�_�o�rb�]]����9���~�K<�E�B�)�A�X��Cp�zO~���a��Qf�!���.; �0	�!l�����r��d�t�1i�x��|j��Lm8|S�no���Xf;�yԭSV[.�n��N�B9�&cѶ�x>Ѷ!�%��!�\���C$�g�6>ھ����Ϛ_�����o/��$����7���wW���-y���G߁H>52�����:��p�k@���s�H����|Y���1][�q>��49?�F���<����E�>k�r	���U����n���8:H6l���fLa�g��X�T�"E�ѳ�}w������^�H_j�'����=5}O���5x���Iʹ]������1�.�U�q>�"�;�9�{��s���I��^.xָ)P;��z�k��?�ͣ��IGfX�f �ߞ�u�&�ת�=�X�"}��#+���Z"�Z�Α?��_'�����pȞc~ӛ��q0Y����Uw�q`����=h���������ϢtD`v��&�_�V�!��b�=�!T,���P��3�}a�>已���2�r�K��Z3��==�]ɫjĐ�h�Mx�8[�HR��H�ʸom
ycZn�\��K~��!D�H{������������l٨k*S��Y_�M������v�z�b�$B�6�Y{�cи�4}Ά>�G���z>�Y���1
f'�y1l&���S�(Z�W�
���T 3���ze0�Ns<�V�S�ʄ(�ZG�F/�q-�n�?��3��Z���F���E����D�J]+���M�w~?=�B}u�����.�ʫ�i���֞Vo]�1Ek�>]���8:��J]_9��Ox����N�j`j��"6�2@�@ET�c]n�2�6Յ��t����ה�]��Hs|�p~)��AK4�Eb�gC;�s��AZLϾ�k�d!��f.Qz������Vl&gDa:��3�Ԉ
���z!#8��Z���A`�BE��4"�g�T�`�M�H&�.X��-Q����p���+o�(0��w�{A�_���𝐗ZPo���
e�W�O;��^���DҶ>��m��I����E&��_;nJ2򦨚�;��C@*�zf��-���n�FX�XƘ�r��3��S����T��@��p8|�(sf���z��	D�Uv���إ5C�NV!E�<���N�KWp�u_����E�R��������L�D�]����m��?#�3��%(�IX�Ԩ炊$�5R>D�A}֢�Ϻf���1���@�!�WY��4E|��o�|!�=��)��t��S�z`�����W�&B���J{V-=^���o���j,Q>5�"7�2�:�M���G�i��13�{	��M�g�36!
W�&	�1?��M��EC�M�V]��o�-�:ߦN"y\�%���z5���;Q+}/qO�����a鈍r���ڗ�מ�Y[͝`m�����3f�.�h&��9
&4��0��|=��BNhZ��͑�r%6c��ׄk .��꯳�W(J���!5[��bꚜJ�e���^X#�jN��س���(�PI�$�� �*(|y�����(Zt���짷RɆ��a����]��y������KB���UX�������1�(m]���;+��8�ߚYK��M9"LP���CB��5d�jh��Z1Ҵ�+�U2�����[����ā�:#�8�.��۰Vʂx7��+�н os��Y9t��r5'��(�����Nӝ���	�����'�%^,^�&e\�?*��Z�ZAU'4\9������1
��E\����'���{x�d��(�Z�z�MA^�v�d����0�F\����M��9S��8��r��aߞ<��$iE��{a"��e2�k��3�QEW�$"��b���_'>�[eT{�Ӯ��J[�<%.#�q�㕊��e�����D����`��>��m�g��Ѽ�T�/ǒ6���Þu�1���=�\1�E[!F��
i��b��Â��p��1w�r��LZ��=�`Ro~�EOzg��DV~�[~89�ð�[?�w��?��|G=���rf�̆W٠D�뾏i�7�R�;�i�O�ܬ�v�E�T��g�mM�Ⱶ�ݷY���CF�`�
D�olw����;�q2x{���hhڟ�^})�:��v��ε�J��ܸV4�8?����qf'ё˅b"#�$�&�Ϋ��n}xK�i�����4b���D�#z��GKV�ۑ?�[.�J�������D`�W^
�;���(L�n�0Ϸ��QK_^�Kg�ː�Qހ�q�N��QP��(��b�'z���n|��>�
�S�y*���!�|@��?AE�\�99_�L9X�o�E��.���������� �W�"c�ꯦda(EF%K�qӣ%�("���v|��ެ1k[z��$���Hm6�p�*�e��&M�	�:�v:���٠����g�P�mg����&��� ���K R��N֧�����G�C�
��l1�H�_�gEUN�lf���Q��F��l��R�7��z�4^��?��<�iòmj�� T�1� z�_A{m�C�Y�D��ؕ��ѩ흞o���SUoKK���Q��=�O�U��k�_�_ 3W��-���<_�o��j�D��vN&��iL=����^ U+�����J�FKd"٪�b�K� �D'(c#���vpE�w
([�E�R}����cw��b�#�j9_��^��� ��)�| �8�����;�yКmn�o�y�9Iagݒ���|��a=g�|w(�"����7f�9��e��g�(5NCF5uz����E���+�Ն'0����^�th]���$
T�.rs��Y�}|rƳGu�iZ��:��wH&r`dT@�� �{�*�ޭ��4���K���[����0-�De��W�KO��h����/���pd�xB���@qmQ����"���	cɶ���p��̮�]���,p��"o��Cߔc�8�~��!d]U�e����]r���� �%OP-�(��EF+0uW*�u�Aw�Y��ހ�yV�U�K�bL��c#�Lhvv��g�P�A�n,Toc,��=}�O)q��k[�U��z��C���OR�/���"UqO^�Ր������t��"��	��/�ʝjʙ�?���-&�͋E�>�s�PZ#��VN�t@��+>:3�WA}�����R�j��{��э�Z�n7������lk�Y�~TrW�!�hɁ��Y2�ZI��-EB2+��н�a��0լ�*+[v������ϷW^hP
�:ޯ�M�Ry31�ꇫ���K��ߜ/���	��Giy��G�A9��U���Mx#p�ڑ�e��Ԯf�G`hg�E�MT�ty߾Q���v(̕i����������~stp;�(��)U�3��'J��1�?�N/�i|��$�>�	(	a),�38�tqᢲ��Q�0�-{N֬ڤ���ݶ�d��h�$%��z���U���jMl��G�"P;gL�l���'xW��~��,G�M�o��T������s٧���$ľ�i�	x����ʝo�¤���Z���o=��e}�<B�i�+�tG}5� =�q�q�K�K�~J�$�%נ�����`��h�4�+����޼�8�˦D�q��7��֤�l��h�~�S���Ay"��P~�n�=���������^ �-��b�f���b�3 �%T�x��S���Y���S B~����/�萔ֺ�U����[(:E����'�(�l��op�O�{�;܏�uǗ��#�`�!_=B�Cv}
�+^5Ƞ_a�*&�o��$��F�~�#@F�����O2�.��x�!hē�F[Gy�6�`#R����y�z�j��=���3I�����x�`��!�r��{���G1���&qB�'4^�6e��Z�#"��W ����Y|Vy�3�� �(�%� 2�*��%z�
�H#�&km��Ƒ��ƭ��[C=T����$�:~bX�Nՙ���^t����})F�cq֤�V����t��d��Hc�(��������4*���>f���g��{�y*_9  e[,hc�h����y�|U#~Ԇ����.�w?9�{�x$�U��Bi<�.����ۗ���O��o�G}���jri���u�}����kd0��P��$^5=��F��|�)4HL���:+d%�����|�D�^�0?�Q�8M�Ng�1D�|Y*a��k����]ƿ�W2�;�8��"s19��~̊�����8��b���^�t�*]��{ˮ:�-\	����%8$�[pw������!8www����������'�`��U5�#�f��S	�lw`�{��8�&�;�̍K�TR�)���:��!��A��<�~DWW)
��Fr��,�e����aE�Ph͒I�d�N/c���O�9C�\fh�'qw�W�!������Y$F��0�0�nD#��S�8����ˁq=ģ�p�ˎ��n6cG`�*\I��ûGsr��O�3x��Π�Y>H_&�I�Z��^]�u�EQۄ��U��,6+�4�Rf�,bأ:6B���ϮҖMfmn^��^BVsI)�(��E0����i�7�K�L��Pӆ��)���\��I�W��3��)핰藦�?{��Ί[ �q	G�A�.ӣ�E#��x@�����̹�ƙ����I���Vy��ϯ%X���V|�h�^��^�b�_c�bNLk��{r�}�x; 6O������^��JHk.Bgj��p���g��:r�g�&)�V
�¾��2�L��v�i�"�	�S#��v8Xnc���������+?��MQ�.�6�(B�R�|��MƆ(�5.s1ws�5�r��0-�fap����,�0�q�����DV�I�����'�KYsY�� L ����R��JC���f�v�|y���u�hE�3�\��27���� e�p�]�W�Qm�bN��8d�MNqf��\#��*H3����r)`����Xrp�΃��D�-����?փ:]h����/���4�jk8M��G��,�iц���A"8�pt����/�!~ز�\Q}���#��h��6|I�fX�T��ۍz�Ѧm�#��؃�<kb���]�LZ�6�,����}�-d�9xk��~ >/sșMP��x�7z"��RN�PF�Ϸ��v6�/nۘ/nM�>���=~��gm�>݈�
�����oue��y�_z���t�O��O�	j4��"�$�?>�Duv#�͈�5%�=�3e��Mͼ���?����wl�Ce�[i-�<�b�"gM�2�6��d�J����>�!ǎ���b�d�I`͂n�]Q��Hvc��k�~JGM*�[�����A������Db�$�j�.s���j1������ʅ�h��2#��&�	���m[���-?�c������k��b
�yl'�4m*.�j�[R�h���i�0��#���:w<�T�Z�Z����hZ��� q�O[�Sh�$b��*V|�?���:�g#H�{�<a��➠@K�����Z� 0�k8l<H|�+Wd��^<��#�0(�u���o�3N:Bšc'��pW���]�mE�bݡ�$V�4��]�k >�t�oB��el�˶��t�n���:9"\�,<1��a�Bk�����E���g.¶:���oӜ.mC�*.��4����a��Kq��J�.]W~��!\��\��ወ�t]?��r-�O�V&e�[��%H��}���CIK����L�Ro�F�����X�G]�'��!c�{hr�f̯,VR�|Y�p�.����|Jv�A����T����ѵ��c����2X�'4�?��D�YR#Agbq^��	ޢ;D�r�G�ó��o������ߝ�h�����~WF8�K�-�܏���ֵ���<�}�C��w�����P��#�]am��E�ݣ�3\|�v1V���� �w6��j�(/kx��aJ����J��W!�Tu�@?ΡQi�%�����	�/�k��^͈^S-a'��S��B��F���x���_O5�u�i	$鈋�6y%��e��2�7��Y��\�ʶR��n����u� ��1E��reE�a;e��8�� �A��_�Z���<:3f*�tT벡'�9�=.S� �ųUY�5��a�ݸ�O�0�K��V���7�`sdw�dÓ!H�'[v���;��9�,�!m�7Y1 ���9Ӝ"�6��M�329pbZl�ISQ���]���d�T����B\�_xTh���y�ah�Ħ:�K��
�{�����B��*�A�#�j]	5������Fꘕ��c�l@%	����|�ɋ{!�R�e+vq����ᔚ�P��-���rM5����"��wn�H��l�r��?	�AC�9}̘k[݅�M@�G;M�=C+2^�YB3\��p�W����C�o{����
/~�ן5�?��!�U�0��/Jm6հ��)��6;���Y�~Ű�ҭ�������I��`B�aH�V�`n������C_+<��"`|f�7`WKt�E��mtX��a�Hh�7��B�l�����J���7�#�RT͓�Pb�b����9C��R�C�fT��Y��lDu�����"�Su�uH_;��]0�y\s9�����ѝ']���gU��#��.�.�"f2-�u��iN�.��e��m���%�oP!G>i�CŘ�5P*����yY��S���sP� $1�lԫvK���W���E�W�-@a���ޭ7��Ђu��ex��h闤~������«٬G��'��Q�ʯ�]�2�ymv#T�=ϧ|�AZ�|��<�����?(ȥБ���o�Z�<��3�و� j���H�e
g�,K٪�w?��l�,C�r�~���hrV�I�/�}wBJ,�A�O��:�Wa��P)�Ϊjʬ/����s�n�1�W�Z���Pl�9�id�C��rײ�����簃k3�@�aK�Κ����q��9� Y�}�o�����~MA�$A�D�֧�E���<5�B����kֳ0��VK�9�	q���?�c��s �hǑ���M5��8�Q5�w��X�d�A��.̮ht
#�����T9?0O��ui�O�6b�?P���>xȊ��7@v�j�~�	癮�%��rհ�Ea�ǮE���tV�k��QkM�DQ�\#����I������N��0��ӏfbQB��K��:h>�ؖ��GD�.�ߋ}o:=����M̕�N����O����]B�9
e/�K���tn�Ω>�818	J����D���v*��?T�
���
��=��V��I��ۏ�_���"���N?&R�ɥjj�+oh�H��/%�{ko��eH�a �@Z���S�	��� m�|�K����ચ?t�U�Wz!6\�I���n6������m@� ��3�~���@�]��} �,2J�/�Q�CklsV/:�O���#�M��j�A!R�(�b�긄.�+�����4��AٌA�g�T�:�.��/��:�~;��{cNmX�F����L'�1���d��|�_���o������2�d�L���0Q�<ʮqqV�c��,8*y�%O	BF37�T��M_x�f*b�4��t҂X�(�����(h�R����;g�ޯ�;��q���g?��@ޔ9R֪^5t3�l �~!&U������HW ���AF�bQ�v.�������ט˻��E�n-xPL��A�j-c��R_
�)H"D�t�XW�@>g�J'_ ���nv�%�yj��2_�bm�L�x��Y�3��^'u<bK��yMvR�!�6�%2��7*���̺=�0�0@�fe�3ďIZǭf�h+t�`gz��X6�E/�ʁNɠe3�-qP�l*����MQ��ӡ)!\��*�����췠�:�O �(7�'`ߏ���\��"5<U����?'=�.N��@�DL+�����"�a���iR�+|�B37�\U���hs@Հ�K����/Z[���`����'�~���c�΃����nӳ
�`�.�1�gT�X�`��p�ǐD���s��I�M�rHD��b^O�a.=kF@�LV���"�wx]����B��wѬO��9�po�N>�ӥ���0h���mUW�2�|���������'߄b~��
RΝ1�?hw��8��߭�acB�D�Ҋ���/�;p�@����\��`��(��07��Y_�b�p�N�q�I��2�V�����0�s:�N$OҠ��`��X~9�o7�A5C%�:�8��]Ed6������s��O+�Y#�����!��^��F��-�S��ķ2�����ͫ<BJn$���H��B�&pz�)�d(6��\�w�Dq����'2���[7�ȢF�3�Y���_~R�%�v�s���-�KG	���m+f�m|}UH����b��[e{%T�u��|ٱ�`�(f��0@�����?���D�V���@�vF��2��ѕ�;v��Xw�޶R ��iުnJ:���F}���\̸=a!�����C�<ҭc�FLʘ���c�1;\4�yjT��r��-� Ϡ�v����7x1U�.G�C;�S��\W)��H��5�:�N��W���
su��G�-�k��Z�9w�[i͡_��y��c����3Y�N��.�%�r��c%���L�I�Me�6P����}��g-jX�t�����m݃^5Q����3J��n����2X)1�t	��r������ј8c��v�޹��l[��h�$����d�����Y[��Ez}��h�ͳ��E���#�s��������r�"�r}n:���!1�m�X����Ǻ��M�ܛ�$_s���"����):������s���wj�=E_��τ_W[�����Bn���� >��t͹=-�ř��~Y �*9Җ)I���?��v���cƶi��E��{�N6�PC��Gi�n�/}��|���w}W�z�g�� �����Ty,�����=�`]\YьE�#���׭����!�tv�uZlT��������ü!�����?� yT�
)vk��}�g� 6���ξRP�||���5�I�e����}zGV��	�ah_�
�J	 ���Z(��ϥ��6FF�ҫ��v�����mW�2���t�t�Y�x4�����%�L��+�a���ٶ�������e�ġb|��w��b�mw�k�{��	tXg�&��d��{g?R7@��g��o�|?<�ξ7����G�&���3woע�,m�s�e�2�?��r#�6�f����$&�[@�P�皤���'�V�X'w�d��*d��f��C�4�j8������:���=�@R=a�����6��������늘��j4���$ �o�֐���S`��ܴu�P0� Sܵ�r�C�x�j�1n͖Ķ[��8p���3s�Bqs$Z�7�ڋ���S�%��Q�i�,糏��7W�qo2��o��S�s����pt��U��#�6�ҡ�����e~�o�ۓZԋ�+��J�� ���zI��Ï��Y��ڰq^ЍQ۲u3�qy�(��cxW� `�.�c�v �w��Ѭ��9|��&ױt��1�[��k���V6{db�I"T�1��^�5����.��Ʋp�/W7��g����������{AQ.��0�Wх����J��[�9p��Oւ@^r
��{K�tN��u�d�����tJGc6��N�G����"L������s�)�0�����2X�+��Q�]����̅�(���!����أ4N[R�����H�	M�c��T
o� �l����z^���\���%+͘۸;Q��{d٘m ^����|��.l�c�syX���Z�m�Р7�v:_مݩ����Y��O�-�rSm��3�� ��s|��X+����4��5�Z[^�س��.CC'��a[9_Tę�'�ݣ& �.%���6�S.��+N�����BC*1-;����1�5�����<M[�2�pzk�h��\ܪ���/����k٪���AzJ�J������+J��4􀤽��¼�E	M��o��˺xa>��/�Nc��u�:{S������t@�{�xr��km��6�ר�{����� �ִ��D0��Z���i�ؓG�8pe=�B�}�@~i)w[����Fi�Z !�i@0�񰼘�`�x�)<�w&~5�ٸuvw��\0�~}���>�ǔ/���(cz�9Kj�ƫ��<#Β�2������w�83�	�oLI���K|�UR��K�5�řG�^:�+07/U!�Ok�� @4��!p���y۶�U=��iM������o�1���9��4Eu��k��s�x���=��|�����S�l��[�PO��7�+�4�By��].)~xn2T�g��ғ���������IZ����iQU)e�T��n���][cv��wxLx�+?}9b��8�篳��o�V���26�����l�DFP���#��lt�������V�7Y9���|M5���B�̎�9�P�yq�:�HZLF�=�@��G�����J��29c���č4F�&{/��Wj؁�����R�6�7O#�y���#x:��$"���y!������j:9
a,�#	�'<�4հtӧ���Cʽ����t+�t-I�]^?Mx-��������1z��@�dP���[y0 �STm���z�����̌%�b��jƳ�n��^��������)�'`/�чO�(7xӯ�?�Z+��v[8��u/�l2�G��Ύ)@�-⮾n����`�;y� �+��{�lވ��v��|��LN��|'YG��Bv�lC�Lۥe���+�r�	��"����g�(�q#�߭3R�����GN�3ǈE�l�-�`�n&�K`�b���K<�b�� ��<	��3z�}�ޫ���d;y�K��!0IC1��W�Q�·,J��iY��a��fo}�|y�?4�x�C��?�S>�'%����M51���g�uG_��7�����.�N���^�7��M?����@�ڝ�K�Q��C9;P|�?,������6�[ߵ���1���s� �:���?��Zӛ��\���U5���eO���d�8GR�v�P_�T-cGΝ��z[-5½1M�^�4��ϊJ h{b��G��
OӾ�K��t+�T1y��sھ�^Q��dءg3���o���������t6"� ��ƅт3��:-Ě���x�c�9Q(k{���?5�3�f��4��3z�o��4�����E�*g��Jc��SM�I���.�E����M
��/�&۬�{�O���-F�]�i��J��᠞ǠDD�?���	p�7؞d�}���?����p:I��ڬ��)K0� #��R��B�#{l3a�gK�Q�((�Ͷ� ��p g�]�)�c�孶%��C��m���E�o�K2��8ڜ�j�<#�[+�U�g�Bd���K!�#kڲ?����J��?���qh�R�<[�Y�X�'� ��^�o��an��W��iI�O�)���v4H�Fm�"U�1���XQ�g�i�[}�R"g&�v&�&yF�
+B��5�q�N��z�2Q��&�6�j�!X�b�#��>Z��:I/�Ą���a��$Gt��$���=�b~���W�ѓ�Km�\�{Ȩ�/#%Au�N�#����,��F�N������P�7|7�v��[ �֚%1~�tg��A��e�rb�������ߎ@��O]MkD�{�"g�M'��7�WtnU���b������$-���-���{
tY@	����Iĩ
��)�a!l���Pw����Md����_4�o��κS�"��̄��-E�N �6�H(�dvP�F[�7�I&ڛ>�kZ'�͡��!F˞�~�	����
��&¤;�����9�[��X�*�z޾q�$ꄔc�p�OZ�t�I�ٖ#@�q�z|M��E]�ifܬ����2O����]� �'$ Xk��� ��%1*��P:��m.��V_Ys[���5�����uM�Ե/ȌJ^=C�BW���He�WIK�����_�l0BҪ��a���,i�\�J��F�j��4[e�S�.�3��Zf%���96k���q��8�H��uk���׼��+�� ���ZE(2vV�(0j�{�)�A�T��HMG��<����l��Ou���V"�����[��G�9	��|��2��(���>�|;+���`�f�˴� ��T�˺ȌT�2�Y��A���EL�h4&�H�������1eU�֬�����uժ��P��Ѥ�J�!A�tT����D��rʬr�st��C�����}Q<|��/�s�X�x� ��4M��G3^Ę�`{��^���ln�'Gϋ��Mܙٖ�,P��b��=U#q�P�r`�M�]�1��v\ U9�@V�~�B%�ǻ���HY����A<OyU#�JU�AN��%ʴ�${���x��6��bq;����	Zs�#��3�	v|8����P����*��|�Rut�7�`:����u�@\j�A��/i��u�;���:e0G3�rl�^?�ж~U6��6$�zj b��a�I�K����%5�.�x��y]`���Vn�9�&�Sw�y2����z��K���Ro�0���8>��^'0�,oC:��6�;����ׄ �J_!�q)K���V?:�6�������/Ǭ1+h ^a]2�x�j����޽���lz��u�-�'`ymL~[!N�ʫ�m.GS��l�JlD�h��>N�h�IYŞ_��=2�nCi�t�p��ݛW�M��P=9?�+y�hL�&b�/����6F�4F�+5�â�t��1)z��c����Kiާ��[�������L^����ӏ	���I�{�a(G����ɷ}��ӝ�Nߔ��nl�3�[ڽnM�L���%�O��d�oݠ���[.�{�4 p',�|��RHF'�]t�P-Ac�����N�V�˰��`F&����G���Mu�AG������N�%%����\ؽ� 0*�#�1{fWA6q��t��K����Rh=����v��-�k�L�,0�џ]��U;��\�N��#Rd�xOv�"�\�G�swᾢ��h}�n�1�f���3����ń�:��E �]����Q4�z���\d�y�~'���X�z�&0뉁<���Ʉ��9��\�����tV]R.�§76\�v��RV5G���i��.��$�BmDiΜ���u�Z<��Y~X�� G��1��d2`6�THv�'���n�<1�\n>�W{�T�� �fW��z��꜄�V2��Y��k����-2*t|И��9�@�]�������Ȧ��<��������ƀ�O�.'r���X��A}��۵����'�g�	^�ps�G���E��T�4#��D�|Y��*���Zw�5�VU���w�2��v�kZI�)w`�]Z�����L�n�*���q�{�I��׷D ���f7��V�-��@?��=�H�*��QY�S��4�k�gMU���=��@ܙ�V��?�PO�Z����8�d���,*C'R���L�1<T9�D	1�dM���1W����Q�y���O�+�f��O2#�U��c��a\�Eυ\6@<�����1��f9}?��%�YJ�,�݀��۞�́��-��Q���4<���RTw�Bn(�c���گ����C��%<ɬȚcc^�*Y�N��%I3��]�&�h�@�W'�+���C%A`���|�|h(>��ܾc}��T��/u��7�̀��.�vus9:Вs{ �IN��Qp�T�rى.���ˆz�f���N?�-���dYme3ۙ�D����p���p:�g�j�Sƀ��,���ه_9��We�k��K���r����*�"�k�ΛH�3, r�f&f�WL��Y�ti���y�Gg&	v�@ny�=�i��A�d2�.�hj�峨A��͡�؉�?]�zvNm�܌�We&�r�SJ�I	sTJPV�YS� �K����Y�ܽ��-s_Jj�P��n�G[��8_8o����y��N�`eF��Q3�ؐj�$���?��16�l�劳���/���!5L�ש�y-xKq�=]� �'�a�!�e���ׂ�f��lsn��r�2	u������2��	=�\�c�)���{_ºO�6�)^ڋ�9> �4�]Q��E��;�!N��D�Z�@��-��wy��UM? n�y�3Xu��!g{���d`���V
L�H�_��`X�߿��W��s��+�"B�X����;ii��,�ו'Sb��d7��W��4�.���ՉR��,�T�)+3�L��ܒn��'l���|��t��?t�V�����K3vbA�����p�7�����YP�B<��PܱX���R[�m��O�;�+���GG��,ﻰ��]�Fky�q��&�ȇj��L�/����տ�;�)հ�����$�B�����X��7b^��@H�\�FP��ro��0F}�7�B6�������ߋ#y���&[/�C���𙐣����3���H��� B�WmV�)8�P�����VI��Rx����75���G$�R��JƩE`��ݜ�ghC}f�S,�/`NAJ9��Vº?������Dј,����E�I#�1Bu�ta/b3���)��������X .�j�� �|~;@�u���&K�u�[_Mk�nfٵ��?'[�� `o�H�,c����f���qc/7�4���_3s���У`�n���멖T��`a���݊`ѩ���"�ܯ��.��9��;m+ʡps=#:H���,u���������$)d,S���� ���B�7��!b&3��5}Q A���h�&��đMsT?��I(�⯫���L��,!X����hʻ���m��Ug����5�ɨ�# �>S� Fo�ҽ^˳�Y�la�M����o�T�dy�)ocM�"Ur��؜���TCz\�,���\����߹1��I������;7(!������2�߹�����܈���wn���������_u�l�0�/T��uҰן �� !�^kK�X ܁e[�Hxǡ���I2~���5M���8�@A�8d��eG8���{��W^c�N�j�tR�z�u ͎�@�<8 
oTd˖[U���{Wn[C�;���$�g�Ʈ �&Or��<�������=���h��s���T��%U�ƜGi5�i|8�?�.�@'�!1�XY�q�(����hX���+�iR��l�0"J�	��<�uT��^�'ԝn�j*�9���2��#y��a�D]�q���Y#|�<�4�$P�d'�mB��|��i6g��A��������Jɀ����|Xyq�f-oBK�j��)C���ąo��Y#�@����˝Ҕ>�]a��� w�tF��O_f��{I��`;������>1���FVH|r�
EK�-)D��+�䳞��w�VJ��CG�}���寀y�Ѷ���5.:���G7�:?j��_j�����_�A��2�&zpl?	�9�F���N��[?�7bҡLh?����5iPÛP�c���n3�#��16�����	�F�]{^���(�֏}����ւ��`JD�A;sL���N�,����6��sw�eM5E�_�m�}�
WR�1����7����z���u(P����ڣ<�W,.c��)��/UǷSQ�������~:�d�|K��F����6p�m�OE}�(����T������
���`H�h��������L�sS�W��+�>�����\���
��l��0ê>b��M"�b6k�e}��M+ҳ�R'ㅜ��F���^����]���n��f P��B$���o¯�oP�"�@ah/����\=t�z�+/�<p�+)�!��y��zȽ�1nn�N6���`��mOR���o�zT�ۿ��C&K٨-Bp�O|�8�ŧPT���^n��ߒ/�4�T�W|�92���yEV'�0�,�q+�т�l�.53�{).��ܖ�'O���>��JO''�8z"�	�k!D�}�~�~'�s�%}�W�T��ߵwst�^{ጣb�k�,u�$an�!M��.I�-KT�Z��W�Ā*����bw�ն�ȝ�����7�w�i|,�������=�A��㌗�7�l̈z�T���;��������Rb���|�8��=z ℡�	�F(�/��H�ЁE��x�?C�������}�D�M&n��=��(���x1��^�B��I^�G\�3|,ݦj��vVh�M)@,�I�+e�"B���c�)�cmP���8���@�P�B��zlݼ��u�+��5P/b�c1M
��l���>���,�d7Bw��ޏ�:�(HKyBm�iݶ{]`�"�i�1�ftN`�,"!�cK.�Ya/wmm:_N��·^M�Ţ���t.�mo�/�V�R�Xa�xQ��4��<�o`�X��������{�9��+m��{�����Ռ
&�nǢ�VxE`���[����tr,M�����c�DE�J0;%�H2�>�t?�x�R���F�.Г�i���q�܉��D�ק�}RL ^x!��)�8p�<<@v�u�� qG�����4S��@}�t_m���
P-��8�D�@y#ý��W3�K��?�f޵�u����5������s6��@%�-!��%*h\�Y���bS�T{ܽ]��O<�{vk*��!���}��^?*0�Л�p���0�y��ye�`N��3��)s���>��2ݱ��=� � f�?�)]�lҷ9��1���j�a�%p���|�̉�F t��<�$�0��r�`r�奷#�$�x�%|��/���ϊ�@�n+<��l���VB�?v��(�6��{���]o���z�������@���?�UqU��<d��M�P���}�I3�Qoݸ��wgs��'Y���e�.�r�ވ�n~���	6C*,Qx�T��i��	c2y�õ�S��s����5������}p�;XJ���}��$v���'M�iқ�4L��PxrZ��j�^h���?�C��!r\�I9�z������2h/��N��L8vj����.,k���џM��Yv�����VԓO����x�|��5�"�=f۷���KV�M��$���[Ž�$yy��i�*T�W�(3���̫�EyAWi��*1F�Z�+��R�D�Z0��žyl�'�z��L*���ڌ��ٶ�`EV+>u�.
;��������g��g������5ȧ[�
ߎ���56l��(��;���mw#�M_��u�*y9��(��2�?�pP<Co��-<�����"��RZ<���F�Ϣ�"�wY�~i��`x��b������X�\�v��ɒ�6�c���µqh�\��{��b_��i{�硾���|� �6�-�f?�.O^-X�6��:��=ZwTP�������bJ�J����ۚ�m�]_�����{Mp���,Y���jAz��G���5/��t�r�Ӗa*u�N�i^�H�Q�?�$�[���H��oկ�p>���+��vxk�Dё�]����/�q���x�r�)���ڬ�KX�`��G�~��7S=<�1�K��0�E�Z�#Du���Ӿ�\²z?��{�=�sNE�f��>���}��eK�!T�);��}����Y]���`J5��e�B��Zq�z-?ΈO[0Tc��ԑӂ}&�פ���7u�Vz����'�&��;��aR4�������Gqֵ穖��sa�x"m��`��IM���`�:�	3�s`z+P��{��̬��˾e��W}oȫ�΅D��j�7%�^J�鮷$cQ��\��^�$,0���C����N���+���;���7����@�na��dUbqt6���>�����8�y���[�h;!�/���?�u�+�"���g�����a�y���Oɾ=�o,��tV��h[+E��`��u���j�L������R� +侖�O^JXOv���#�>���~(��켆��_������g�}�]���.��g��`s�W*ݬ&�+�t���cZ��+Id��x��ހ�@C�V�E�Z��a�I�%���o�N��)�MR��@��)ijIXV��J�h��~�ΦM�����2�ݮ:��8�/�7K���ܟJ��=�2����[���a	��;�5m��5-��QWj�R��d�O�1
z��DD_�B�.��貸��8}q����&4��}T*���=kj~�q��|�+3W%`�<s���ߜ�T�r�d�'>l_��� 5�gSP�X���u�	�`z��J:4�*���,�T�5m�6m;eu�F���P�8�*d.�ꦠG����K ��D�fmO�lP��r]�&e���]^��	C�l���y�`Q��4����N�M�s��2��S32����k�b�7㖩Z�V�=5����~�ߴ�>����5c�ewc[�6y���D)��,��O!�v�Ijso�ᦸ��Dj1:q�3�d(w��.���W��RX^�ws����on�hvT�}�xG�q�S�ě�C{{J��!ώod�a��D�>��g,#Eݝh��sQ�fj��E��V{�k�N�"hp�A�#JW���2a�ba?�lj�b��R�5h��{�O�oǁAwEFWQ��8��8�_w��'��$�ww��A��;���r���bB���<]oIxi+lv�%}=�e�,ҚN;n�j��_�L�d�"���������U�����+怖���'̸�w;��6#@�\���I�[��5��P�%3$/������w4��s
��
��x�~�h(�͢@՞`�T'���<���pnI ��Pl`'+'�� ���XӶ�[F�֍wفO�|ʠ��+���q؃��%�ٍ]�����̏&a���o1c�ɐ�����T�/��ο�D�d¡�(�3؋��s!w�B�6͘{F��&O<��[Y�w�F<$�ME|�5�ۿ��Q�5M!L��зLL2~��b+i���Z��hR�?�t
�+�{;�w��͎��m��@����/U1G;�'�

ll[^G��?��N_z����±���|aCg��a��j�x�Z��x��n�+��|e#=Q�i^y�k�8M/[Zǆ��6���B<�A��i�7;n�z?�y��������X[��ʡ����_F�lnv���$�i���~,��hw�sN�e�m������۶�allû��"S��f���F�ҧWa̷���X�����r'%�O�����r���|G�Sґ��n����HW,�w��N����i�QI�!�q�u��F��o	�h�'�n���oEu>A��/r蹲`��p��BB��6A'X���m}�����B.���Ħ�eC��W�Er��y~��#��iW
�&| +���ڵ#�gg��;��M���v2�:<�ܳM���4w:ԋ5���g��Ev�����Ք�I�:��m�h*N�:M���D-��E���FW�W'���t�u�/�j�D�=Wc�!�Q�x��%u����E�JBk�"��V��S*@B���I|M��?�0m�5vHn���cM�I�$P�& �9�C��N����*	�[j�%g�yUj8��6a�L?�T\�u7��\���T�'ޖ�h{�r�4)�lZh�*�uu擓�����l���C�}���X�w�9I��ON."���h[Ph�	)��Q�LL�����,���7-| ���9��-�c��?���l�����},$>v��z6�F0s�`p��(���Bt�~	&�U�#-�BS$t�Z���u�#ôɴ��{]�PF�Ta-BO��` �ˑR59̬�Z� � �6+��S�ֈ����tT��[����ޠ�0:�Ԁ�����$w�a������©f�������"I.�T��\����Q�oz�&����{��1���|`��^�1$�u��f�)��<�� /jܳ{�k�U`�D_c�&F/̧�,ȁ����a��k���ڡ�x��o���'Ɛ�C`6���\%���0��6
>I��ܾ�'ro��Ro��	���U�F��jf�&��JC��ow��h�u[W�)G�0ub<�U<������!����ٸɌ|dW��5\S�۲�^(� �(I�P?1=p���'oC��u�C�/�Ƭs��Kk�{��b�`E�;�H�(����s��\�a:�r�[j�!��	��O�� ��s�rd�c�%*dݒ.��8�Z�Rk3���v������1��~�_�_��+U�7
d���2p��?Pt���'��Hwu	�L�3������7A�Gk45��ߞ���=5�$���_�]�!���b5����Fn\��n�0�<r����˹'Le��տ��9��B3���%m<�^ly�,8���om�ʔ.��0��x3vh��r�E"8�yY�/���0��S\�����n�8UM�v�9��~|��M�JT��t�uB���uS�S�IB����������8���~��S�9{�Cͫ�P'��##�]1�
�P1z���x��iiq���񆼠S��D+gR-�Iƈ�qơJ�7��c�O>����}���咥x6*����!��A�b��k�H�F���N�����u��(za�%�>���(�PcñZ��F����^��QJ[?�ZY��)� �y�����^CL�iW��Z2 <x�_�;ip���&˸x�>u��Gp&Ņ!����d�O�mgr�l�VK�yv���E8�:��sV�+cu1�?�{���$���D�9o��v�e���q�פ�񐨵�&�nl����D������+��A���v<���0���Sf�������Y n�'V^J>Ā#�~�N�Mu��<�@��i��s��{���]�*�V4�����E�F�I�y�� ���� (�b"a`H�,���GN�n�
�jcG���ĨbHoV[Qf$��*n�4��r��U>�LJ�m0��P�����S2#C`ڙP`J�r���[m��t�"�x�.1I��`/7˘�Y����
�F��Ep^�lf��Y��������99Z(����2u�e�CI���7�&KSG���HM��|rz�~���(\�w�#6t*�r�����6=�	awv9�0�$x{�#0x�o��>�����M�����I����G��kb��D�oH��eC:�v���(l����E�jf�H�`=����������%���D:7�  HwHww�t�4�H7HK�4Hæ��E����s����wv�5�\�y���\$�%��I�h�7�]�"�Ux�.P�>�wB��ľ�5l�禯���{<�mm�*K@��B�2B%�DBJ��B6ڨ,~j��u�� 1��(&��h 7'�/E�z�o�K�S�#j\D'%��
n��$���]�~�]��$T����Jo7�eޙn-���a�h�L2|{�Mo���K�7y=��o���{��<w����F���)$(���<��}�*U >$��ޣ��M��s�	kk����'�M� �{�����S��V_��c���CaZpZ"��]���#>�@����;�jbrK	�j�cCڿ)���xoF����� �pM��o-����v��Dk� +b��T���X���Ѻ-��s_��Ӗ� �K�����+�����.)Of�\:�.�}/�����8�g��c������0��w��8���L�Q�)f��>��¨��!`�7�6�I_ h3�4Y��CQ3�SZ�Lɏ/m
!�����4��Y��(/l>6	4�+���\&�N�G�����4�q��Z]��Ӎ=�Ў�����-,�ZA<����9y��G��Vo���+v����02�Zv���v	��5�\$��ڼ�a_Wx�>���Ks׷,�ήm����zyzB�B���-�XLG�cߖ���^�4��R��Zj�NM�tj�uK����d�@�C#GlL�s����	 � �Ԟ�f����>���6���a�����h�wu��~P , ���v_+�"ۄ/�\y�_��XH�f���m���M�@ʂ�n_i���%"����H��	�ay	,���g��'u�O�ɍwr�pĶ�W.Uh2�?⃌���WE�e,�;����e��JR����,���nxoP8�p�$s�;�F��44Y�k#:�>ַ-��%��'Vo>
��˭�"by��� �S��������p�Ȅ��sg����F��Iv�'�=��mS18�xG��h�y�W�������eB`�z��D&g7���Z�CQD>�ű��������P��b��qjg]#u���i�����ō��d�"������>^Fk�����D4Oƥ�Ҽt��Y�.v��Ƴ�I�<�B�>חV����Հ��7&��޼95���l���	m^gީ��l&��`;:t��5q���$��@	�����,����M�����_���5��XV� ��'>�޸���}M��??�؞l>R��]#ML��NWf���� 4H��+Y>�������Y�]����ڕ��4�-Mv��X5`�1jր���I���(| ^rܩ�I0���aP�4�+O��Y��geˎ�b|u��|;q}�����!����I�z!q���4�rbo_礊���1t���e�+PKtƼ��:‰s*R�\���ҤM�	�Ep���1f8 �������U��A#��%�{eQ�.ޔ�r��!)��
~}E�w�`nͥ��dt������,�'��k�O��-�MY=���y�y�7t��Xk�P�vpm~:bc���8�����ā�j�1��N���5P�j�]�������w!"�@'�o7��4�_����E�6��E2xE%�7[� ha�|��=^��S=?�ƺ~��Ex(��9#�X���0�m��	������{Е$�~Ǎ�m���+���~Q�W��ހ1(�τ�q�5�t���z�t�� ���ǾlP�Q���7��ڋG�N��xN������V�����o�	�P�흍�{d.�L5p̿����Y���%�t���J
��p�IU�juBC��X��;��׮{��A�9!�0Gޑ]�\P�O�?��4�)sG��~f�!R������X�o�8�(Q�g�Ƶ��-�	F'�z_���G.��T�Q5'������A��sC������3�H^��+[�Z�;��DˬP%:�W{8N�h��m��� ���½�%e�:�OhaJ+���[��j����.a�"H������:2���6�l���� 	��6�k�sQk�Q�++��{*�{���G<��N���o�̂e{yW7@4r��Q��P�-C=�OW^-�f(��W�%��f����K؆��z<K�M���L�s{=ن� '���7�SE&�w�����������L���]M��@�����,�%fB����<�/R��$t��b�kQӨX X���渞��u}NG�	le��+������/�ǋg�I^�+]�{�A#a믲x�׿��:1��,Q�=Ձ�tCK*(b��s�w~��Ý�w�k�o�R�7*�/��\!�1�ݸH�d�^�VS�=v�m��j9���C�RE�Oϩ�w�K?p���"�]{B��HHO��J�.���o,�o'�͟���ӣY�?�f8��`d�x*�b�3��*JAr�_h�a
!�Ft ������)��\Jz����/"� ��D�7��z��2��*Ʃ�"�����KV/�s��(}�6��9Ԩ�r8�CԵ�^��8y�?v���(��W4�1Cl�R���W�U�.��)ó
_=;�z�5u��&M�ߚY6C[�2#����У�#?,���#�5(��H4��?��l���c4o��B���ǎ�R6�4�h2KJ��K�3'�:�r�LZFG�f�5�1Y��]:�-g=�%��3O!>���`:)8��[�N*��S�rc�$MVg^Wm$���C�mf��1��,�e��A���a�
X�-ѫm��^�Aa��eQ�a��k��( ��ݜ���dd��P[�j�bþ�y��m��
_��z ��������*�yQ�(�d���w�M���t,��Qk���e�B��7%��M�K����'�xȯ���;5�����+�m����FCѡ�ߓ������������w�pފ�F�%&	��C�O��.xە��o�O�	}@��f�%�hU:�pc���=o2�!ܛ{���!ʷ�"���w.ho�=KkO�|�|&����ݭ@r������ux���hF���x��V�'C���������Z�}L�=4-ʑǺ���Ĉ�ţ�lZ�,<�y���E/��6��ߓk�v�O:V��]������E���w�Ɗ��f'�*B��q�����AA��������N�$R]��W�H-�4K���� 4.:���5s�iu�#�}d�[@	
wv�s���^�u�_�4�T�L��L��Q���p��;j��*O�U;����͢NU�ӕ���c;�w�'�Ӫ����H��F�L�:Y�;3VC�l1�S�3��	"p��s��]mտ�����n�9�(A����K�8b��U%�@M �:��<RV�ni.����z�xGڥj^�P�I����S��3��~�����I��asFX�V��~��	&|Y�p;%��=%��,�14��,�9����=�K��%��ݏy�~�]n7mF�Աσ3�R�)󎀤]��q�e	��io�|���R7�?���x��e�W��(<�.��Smģz�E �q�׳��/@�˳b�
�`�N��b���Q)�Ӹq�35�;2��%.ⴰ�KGw6��[���i�Yɻ�,����5
�7��������	�J�h\ 
���
��~|qWgLS=%��aGpޔ�H}�<��`�Pa�u����� ΀�%�M�� Q���W<��˨�*�.K%K�;��3��ǫ
�^%h����lEy%6��������c�m�-�-��|��2���=�(e��bze� Uh"�ɸ��`����9l�0�\og1g_�
V�Q���ƫ�
?�x<�sk�������>Bo�\��A};J���&�%d��a ���o�ZJ��̐|3`���_��t�`�]�~����7e��ҵ��g�.�̇��'o�� �����́p>*�$H�0no�F1���(�!�Lq��|�YN��Fsg�����2ٲ��+��$eJ�%�_gߥ"Q��A���\�n�u�"�?�L�z�T،;Пg?�8d'(0�q�\g�3��>��p�tS���\�Zr���B��d'��>~�X7��5�����e�Ƴ|UOO��f�/,��M[`����S��̡���g3QS������'����T�@3�L�<F�*�}'<����5Z���y�=��K�w>�E�$q@Nն$e�^��y��B[�M_i/ᣒ<3�Rk���l{�3^���L�q�NS3 ����v�^�{U��D_�����Iy��@_�p~���ql8��E%�.���g����ī�n@�d�'{�iou��5(}�Ӳ�qQ�
�j���'�W�'���1���M/�x[o=vL)�T8����er%/�|G� Df���;�,�&k�%k�o�ɭ�,<��&���K9����;��Рs�����D��T���R���U��B�(���>i���(��'S�l�Y~F�զA�hZ��So�k�&����ˋ���M��*�� É���,h���d�ڰ������GuJ�.?�eb3*��mo��(YZN�����v&2Q��c,��j��>\���;�%�h��J�ׇ<�������y�������tlD�'[�v��6q� ��(R������[�qa�h�m=8*�����f�fi�N�i��0o�]#HH�仃���'�/�~���f�h��;��S����c�m_ݺPb�oM-�����#e��D��p�M��ֽu�>m̫	�3l�}?;�w*����v>, ������m
�#TӲwkX��M�u�i/��!�׈io!T�D ^8��S�sP�V�q��i�]�xFܬ�D�~��Ԟ�tjR|���B��b 0������(yq�e;�T� ���i<v�����4�3z$zʋ�[�������J6��Da�	$m-PV��i���Vn�ܧ���' �D[Tfw�e��{���m�H��v��-Iv��2&�����VJ!nZD�����A�xP�c1��,�^*lu�����s�U�F�p?��N"��?\r���jG�^��A�=���ǞeV�8�5�\F �U���{ݚ9�m��ԓg��"�6_�bpR��w�ߐ�J /C�_R�1�Y��j���-��zݗ�pA�*
s�Z�y�-l	�.�Y�U���iLȃLr_�y�z�w�����+>���R-��̝�)Q,Y`O�#��aج���}��+C�W,�	gvK{�L��]c��y�c$o�BGP ���I�ruo��`���MI�a;��s�ʩ�v˥[]`NwDP�Й���}MfH����8�\���n��"aV�+�ح��S�������qt�	�^��I��sH)~�\8��Һ��`��:���u�a���)`�j��eV.�p�w�D�T`��w-Jfv�N���=}h#Kn�Y�W ��N����L�ߓ�N�9\�=B��d���B�z�Txxh(!̑'78=/˸;���<fW�v�-gg-���wz����y-͡�f	�n��"V:��R5\��F��F�M����\,_ݖ���ܽI�S)���;��U�?oaI;�8�ZB�&M�C���Ж��5:Ya������9E�Հm�66]�\`�y�w<H�+5P���h	@�a�Z��9����y�����|�K��[3���ډ�b��A��Z�X��+�ǩ�׾��kL�L�T�TkGB���j8
�
�6~���G�����p����M�d�/�h±����!�����St�jp�Q@��B���ͦ�e�d�&��&̳�
�Ύ��I��.���~5{�=�bj`"U�S�g����Bd`Ok���	@g;��W=j�!^P�Ӆ��zJ>zA*�s�� K0ֿ� �*������Xn`���;�b Z׉c{�ĸ@�4z��<���c�E��-�J{�(CǠ��+�F��\=?�2�+u�!�	#�VO�(�	L�tNf��q�r�z�	�=�<+���6�~� ���~@�8A2��;]c��x�@T�;��Vn���Ը���K�20nt 
Fn����ElN��6@����L� ����/��]�(�!⍱1��O�����{��V���da����%��"�����Q @!ʿ������|��t��ovD����~����V�g�X�+��B�\����<�t�vK�mq�m���[�rVn�����	.�`9x�������{��:�+�t�,*L��/o��;��`��)�������!|��HF������h�HO�Nƨ i=�97����nwڸ��leGMv�ۊ,Z�f��#CjE���.|먓\H���@���߉[��i��ks1A�TZ%P�����'y۫>�v�^���_2v;�ة	���]���6��⤥=�|Cc�7:m�\��~�#�m*��CJ��>���}iI� j�Ga`;^�?�%�L��D`�W1�wƁ�%�DH|��vަ� Z�@,�HB=�����3�����w��Qh���1w7n�gN�C���s�c�z�n��Ф��]��H�}}�o���⿜�� �3��,��)cL:���_�Z�V���]!	�����C�.#��l��p����v�ү9I�ؓC�F�_E;ʍ_�툈�~OdH�p	�*�"2)	Kg�/����&~�[h�̠K�A���m��_H�]�s��`�;.<vs�&�7�^�g�L�qȕ��	;�-�<'A�{��緜�u����0U�Q@_���R�;�az��c4X}�:��Ii���j""*��.ˈp�[ߍӈ?hԐC�W���Y�Z6r��}^�b�����V]�Wo��l��D���=Mځ_ӥF��'dmN��7%���E���7����L&"�~�ژ��}��瓉d� ���m����fK�9�<pߕ��*<K/��M 5Y�4A�����%��	���d���s��?�6$)ޮ��3�-�)/2�{�荐KxZ��~8�Y���!x:l�8!3.ی^�<�5�'^�W	M��+S&�ѡ���Y�@M���M�Vj���w�'��<�i�4���oq��Z�ԑ�z�4�L�a�ϖ����W;�d�۱B{�Aap~F��(��1�"�o�kΆ�X
Ӟ��\PW�y����2���4̿�
"1�ʔ� Dl��&��&��
�w�h-�ur�(_8P6Xj3�l���D����(�d-=�C�((B{��PB*���-M� k��M>��a������ǡ��Dl�d/�0�������m�qt?8�pȏ�.9�Ҡ���[r�aptc���󺡡������n"��EBW]�)�X�ge2>@�6�^`���Qo�o8^����Sq8d�vIӣ?���޴��"*صG8��-o�����ʬj#ЃP���*�l
��(F�k�5�S% ?�p�郌/8�Q��I����+��� �N��m�ݤ��4�ى`�ӈL��ڡ�I��H(��k��Y�0����	�Tu�Xd��,��ڿi@����w��ی��/�͑K��z��Y��F?������J-��_�T��[�%�z�0��V<B�\B�ȩ��o�%��Wlg�����c���$!���%Pi2Ns�  �b��dsXA���|�h�U�i ҮX�Ww���
�o�Bj���s���56K]/�վ~^i$?���S���d��7ʶ�Ksj�r���.�L��2F�7�	�P�z�f)��<���S�Nw��ڔܐ��\��_=W������Z�Ƽ���:�b����]B�YD�w��qP������2�>I
ă[wjEuv��휱2��Cr8�RI��G��� A���o9��ԄL�&=n٧3ZSǎ+ec� ��97;���L	��5��7U�5���2Su�c+�i�dg��xT?6��QU%�Hz����8|;��\ւ���\V�hJ>��'��$�-v��d� �NtMR�m�l,		N�����D�a��R<%��M&���*���c��9�ENz2�c�JD8X�]�G\�ޝ����X�L}kbH����&�ϝP}+-��yhJ���u::�
~
���Ú jf��6�e�@�EN����A�cS�Q�8�ߦ���d���14Tk���ݺ��%�Qt%X6v�M-^�YC���$Fx�H�DH�|N��[~����"|+1^�}2��2aJ��`/p˱�vr��>���(3�&���G�m�0]��l�s(�䰢�R���)�qq��J
Gj��љ?!�^X�7R�k-�⹳�ԵS��$��#ލ��|�%";y�����������?�׿�g�\����Qw7�ڪ�e�����硅��5���^f�~��ً��GI������.c�R��G�㻇C��d��%���][RH����
a_�$�;)Q�v�]u��{����ONWww��P�����L*'h:��@���kV�ܞ[^�������jZ�y0L8�bş?���t�k�uh��!v�F\�oڭ7@C�FHJ7�6Oj�U��9@�;��K�gw�b�o�#3�s��rv��B"�./R�d�'��m��T�qE%�����n��J��k3d����:���7�|8m�|�?4�L}|;v�yW�bq��1�v���ţ����A���W��"�L��xJ�h��^��{=L
�o==<	c�����\�-���n��-���z�-*H�6[�~��e������Ei�F��0����՚1�����*ע�x&���/�,I��b��K�$�v��g�I.m���g���^�x
���S�Jî;��@$��lݴIzJ��O{�o�ʾ)�S�j���K�K�eǁ���ʓ��T-�>8�;���w�jZX����:���S��'��R=��ے��l"v ����kG��� �n��>����u�feH���g�H�O{z��2R��8L��ct����GL�V ��S�u��7��n3���X^M���e�"����E[���\�/"�ɯ���8�U	J�ܬ�r��D�F����_Tm/N��'�N��0����a��K����1Y���*U�eEG�f����T���^��'GP`�;x!�\��ق�Ηa҄ E�"U��j���X�O]�x��$[�(y�Y�VQ�p�G[��F�2�&���D8��0�/"�˸ 't[���	a��A�pO��'B��!$P`2/�/���/ڸ~�m�rO�������?S�9�YA���w��2D}�]E�Ǟ�N�/�`��P���߈��יƉf���o�Zn�����[���C1�;Ǵ4;�w�5'|�x��0�	�q��t�אZ=}Q�d�O޲+J ��J�Yt������K��{89�<x�#{��Bb3�ޟV}�B`OQB�L�:!J�<p����q�*���yP禿�����㊈���,ٟ�����,�9�t`{J)��J�6s�R�a������,t'����XX?T�������Sa=Œ��|��O*���r�Kڃ��L�s��$L���8�s���n���ξ�h���{�K�� ��܄=���y�z�|�z�Ք�p"|f���D6��(ͫ�q����k}����4����bu���~-�]����0�J�95ԄF}1�D���#q��W�~1�jl��l[!*ʟbӢ	��=?� %�[�����M��V���Wb�w����%��n/v�J.��*ʹ��BW��Kpߡn젡�L���S�nD�A��CV ��r}C$?��+EEvR�s�zr������u¿��	�i�̲&xU��o���L���:*�OQ%�d���U�h	=���s��A`߾>;���.eʱS�0�k�Lߪ>[2�z���"� 
�f}�����,?���ɴ?��0qLih��x��#mP�T��ߋi-�/H�K O�>��2�M��X�wmI��<���x��V�y�Ew?ʹD���	���T�l���<�銺�C�osG�^�I�Uxrl��\�4;7Qw�F��b��#�VEFfm�;q`�J�}G�6�c�O- OD�0�k�Z���8�gj��D�gHk�Rڏ#ΤK�:���W��~�m�\�S��2\�%�
��.���S�؜����0It&�������G�d��U�ҋ�9 �']�������o�"���;�cC���j4H-���������S�̵��c;v�H���ٳ�t^	��T��g������'V�	{����RT���GB�]��ؘˁ)9�b���E��-���,���ɷپ�Q�$���b�}L&[~�f�q��ůY�z�]O����X�K2Κ��R"͞s9�����n�h���{J��k�4��	��a���3��(?���?��6w-5�s?`��}(��n����;b�}���a�#��^z�XC��#��e�ϫ;Z��;4Y�nZ����MoH��֮ݭ��
-�EmW(Dn*Q?�<�j ����L�]dހ$rz���T����h)ϋU��1��K������h�.x��~�d���Ĵ&�*��x*�� ]����X� ��|��_ɶ�3�yxv'�byV�aI1���8������n�|gm����x��N��BsϠ�}�٧ �7�ς���'�D�����y�����|�7��	ۿ<��0��>�^	��<����;�R�,U���O�\[yvdaJ�6P������)��jL�G1�o(b�.��+�6��AY._uS B7��ċOfs�E�Wp��E��=�-IEKJ�hAe޻�1�OYH���@��bJ�t��S�c�U��DiC{�`5ЄW����>sěT*�9$��o�J���P�rdj���(˸{L$�A=ޔ;ȳ5���;��@ʯl>R���R�~��v� ضϟlzY)|}��peM?�g�5l�H8C=�R��3o!?�3��/LH*+
� ©C�w��n��IF�S�/;�\���w)�5�T����?��?t���s8$"m�D#�ea:��p���(F�O-�8���"K%�;�x̘�h���� �X���R�=p�T�W��s%�Q�9wm��7�L&
c�'7�4���>���r��Z1�����2�y���X��.���+|?j�"�\��έ���d8�&}��})��``�^$�5<FjKوs�w�����ˋ�r�ͦ[0�<^{��-�OZ}�gdy���x����0JQ+:Gt&D��, �n�ݾL�lz��}�b�0�9�C����J��{qlkY���]��XvW̩�޾E�\�쑧~��Vw��Q��P�b�� g�q�/��!��	XĈ��?�O#l��,7i���_�\ ��0���Q�h��;���hZg�e��$��6��]�Z@z��f�i�Ov�M9�7B���%��js�Z�o��n|�>���c��~ӯ�:i2f1��'C�ܜ%$����%�z\�EC��~Cᰁc5�������X<Y퍔�(��Ҡ�p�I�=�ו:b����	����E<�#��[�-�p�3>�Sw;Rg��*���u�"u[HK$�A�����oF`+S�1~�ʢ@*��2Ka���j�L)�2�Ct�*'nPM|��X�H�����V�/b��$�6���Ǝ�!P���J��h�i$��͢��H)`�a���a�_�Z֑��.I �C������Ú��mdlrJ��:�z���94�m��������Aȩ����gă��v�ϋ�N�i�j�D:S" ���*��P�ң1�30�cO��Dr���U�#��t6k(Rubd�r}�ĸ�v��17�a�
5]~��$��c�74��}�y.�eݑ�}����A�G,V�+���et?#�뗤��֓&� ���>+a'b��6�P�>�lc[�*�W;��[@N4`��?���� �2Q�ݗ�_�9�R(Ͱ=�Ő�V����_�o�)��J��	�o���h&gn!����=������6gkV��1W14��^Ox�(O湺�C\��7��k���f�����̩Ek�+�@Ye��1�F��	�+��G1D�@��0�!�K��[���;������}�F@Zl����Y+������e��]���l�q�6K�f��,R��v��*���E)
�e��:�ܙ�ά?_h!�\-D%�HZ���?o��� �	���,/��AT��EF��D=�:��T���,�z6~��RxưE�P����e6�kNKɇ�[.2�{n��\���噌��sj6-�������]3O6�E]�ų��T���,��a�|i����ИMQ����ןdɔ����Q�MR����l/?[��r��E�����ȑ���cL=��*�`fɳ2���۬Q&/����O5dqE��}��m��=���5	H�����l~�x�)��):�q���0��~G˱釻����A�'����|H�>�U�Q׉+/-$ ����^�%؋y9[�׃�z-�5��R�����p �gix*� ���m�Z��
���nӥ�Ryb;�Q[��F@q�5l���~�ō��UH�nw�����~5���4��-��^UJ}�Vx;U����s'�oT'��Q���b}D��!�@���^�X�9�c����uQ����!姊���h�������j���k�c\�7�N�G%�.�O	+���|���bg���k�F����3���\5O��=�协_g�V����h����[��-�0b�9`�i�S}w��{w䈿.D�*�	l&�|�2�P������h�w��7��&'$طN�ڰ�ն;���w�1(�󔎩sI�\�PO�f�G4lrDgAZ�!���o2�<�;7{���ݮc/iGU�޻Ė�=�r���բ�/�ۺH:wJ���	P�h�sk�� e��:Fg���	����+�� J҅�e8���i������������ 8�U
1K75��Gt��Oi��K8����^�cR&�K��)�mI��py��#ꗫ[�*�H�y����f\�����Fl{��2|�i- �$@�]T��^�/�d]F��gޡ�h�~_9I�ǥ�����~� �߾kY�i�jȖ�-^rD��T,��#A�E{��/JC��}4%:�©�w�ϡȐ��5�Q��|;[g�6d|������>���c���k���6�.a�j���+o�
g)vғi2x0.i_��09����iM���·㚩�*;�ܞ��{���"'>FA���ߣ-~��櫦��OC����q2��}�B����4�f˭}~�Wvi2e���l8H-����Iu�=�� �W8��p�M˸4K�x��vH�pY�����ޘ�oAJ'J6��*����)��!��W!���KԲ[޶��e�[p+��o���A:�줪�-�;��HO������&�I�s�{��ubZ��/�
WcP\�v
a��#)�?���X-���^�-����F�'y�O���{#��8*�l��PA:�v_6��>�r�l̬5��g=����jk�@����W	�7�
��~�")x͂���pڭ8�BM0\3j�� N!�E�H�Z��L�������p�tɷ��*�7�	�.��)���ƒ'�}���!(r��2.��E[`�h�*H4ʬտT��z�Й������v��P�B˯��t��t��d!�G,0*M
���ܐs��{�fEkίc��Y5(���ȣ�zﾭP�$Slr��"&�9w��҃i��A�~���>�6���Q|�tƚ ñL��V$�0ZGriy9zL����z�l?��X�*��H�?�&���LE�3��]\k�b�(���e[/�����4�O� d3	!��d}��[�"=~�ʳr�c�1��=��\]��Yo�fō����~��	�NAAj�"�VǫV9�����>c�\?V4q5��u�q�\��y:�>\i�;6a!c��K���������Cha�R�K�Μ��
5��)�Rovvz�emj#��)x����U|�i�ʖ6��od 0h���L�4c=4��i[�w)(_]..5r�H�/�a��p���\Ѯ�HU�I?���&.>�$�a(��
@0����C����	�?���*�������w��}�����G����}` �
�G
_O2���&���#��N����I�Y�u~��������q7������o��R9��Zr\>��=1��ds��
uw��n��U�$�s��v���:M����NS
���D6����4����:M�@���N�}���,�����4q{B��������K��_JxL�����`�l((���겪r	�6"���əި�6�w��t��2[�V;q��p��<Kh9X?wP�Z^"�l���Vۼ�O��s���U���a��e��	[��gde3�5OA���ZK������������"��Z�y�-뷝d��I�z�
	��r�R4@е���\mas��?d/֕F��ow^�|�uU�0z�wc�����gI�X�V�l��f�A#�=�)1V�h]�v�D4�CN#>22�����7�{�!��[ג�ת�*	Q]�Gq<3�v{��^�D[{~��ީD������\��K�6�u���$��r^�r��x��?�O��w	��>�Jm��屣Z�L,Z37F�@�9b���(,Y�~L�)������+r��m󒠼e��UVp��j����>x�\��T����i��ɍIH�/��AC�сZ_W�~��dC�r�.+�?o2�j�Y���a�S:N��Vv�
����4�����N?�0y=0�u֚�$[|e���(H����������kIs�2}5�
|iBx��"zyڏ�B'��e�d��a�jw�{���UF���߂�����{4O.����7o�,���?T�4�"�C�ߑ��Ȧx�i�q��/�>���e��H�1�YK���4�j��0�H�*�k��
?�1-�棼�"UeI���
W�paӹ�'x��p�Ǣ�0��և��_�~�J}Q'�x*8�������8��v��m~'y�3!R��G�v����7���(�[[���g��\UJ�o����H.�Hh�t�ֻ4�:L����?I�P���Y���.(`���R����f�
/?{v�K��%��Dl�>�xG.%�n|�#*�I�g�7l��Y�h1vE��Q���p3B�:����f$����k`�$������}�3�\|��]���k�B?�z�&�7Bj�si�¯�u7Bv(0>nM��Ʀ��5��%��߃$��o�����#��e!yF\ߖ7��cћ��?��9O`�����,�,[g~+E�����)����H�p�K�hՍ6��&��h?��|e.�b|�-ɿ��0����D���k��v�����~*���q�� R-x&b�GAX<�B�A��������BB����O��j�a���v��tg�w@Z�Z¥F,�1)��G�Jg��g�Ļ��KO��	x$?��8zR�����t֒�×��P](tqٰ�~VӬZ�V~��-����{���G4�ԋ����,��n~��Bo��N���0'Զ������̑�0���f��
�I������m[y�+�nk��[��|5�#q�;�MhK{��d$�9^����ꔠt>vl��'D�^�.�~�8F�	�[
����$��KQ��K&C�̚L��ɶq?h����ߙ���'#D;��8����{bcP�ڔ�C-��ߪn5Bj��}�W�69l���|�smso|ʡ��y�`�\�m���#��ߥ����F~�^��+Cbؘ�Sa����=��ժ�ZӲU:�p[E�#���ں�>��cģܾ�1�|�VMwE0��ޗ]���zO���0�1� �zu���6�~�NL��E���;M݁���[��-�����=YP	oKރ_�eԙ��{�����m�r�WFN���A(�U �Dhv� v��4��3ըƪ�������`�ԙ�{�������=�� ���������]��o�vtNMz��_�H~�P� (p���[?��{��� �:�!%�����h�)��V	���8�3΁I\�Q�]tC�iyc<�d��-�@����I�����ģ���_����[��"�V��J�Π�b(X���b'��NP%�ayW|/mj�,�tx����VTg5t�48�W�C1�
5,���r��O��B�z�0� �}@�1~������	E��b-�n�'rxT�Z��S�����}aE����8�J�h7�n��T�s�`j�t��N,B�Q�����T�SQ?WR���_�ު�XQ(�r�ZF�_��������έ�L:����1T=?i��M]d�\{IO4���-ڹD;D�v�	���z��u�-}��+�;�=q6�H�0���ߪ��t��!����V�\~-�Pگ7<A��u���
EBlt�'!��/{���}j�2õ,y����42�q;d�q)��� �.8�\<���E�r�	���t~��ZN,�nK��`{xd�Ў�ޭo&��8�L��v��Hy����������?$����n�~2N��V4#a��߾��?l�k�����L��4�n��r��8�&���0 _�N�S��
[�f,����ҺqF�&��D���(��&S�KD16�u0��	/&|�#0@zj���}�s�p��ϙ�FdM�s��Ê�j���6��,�_�g���O���v�*���z��)�y豁����=�-mFx�	{��@V*�	�@����~A8��{N���w9���x�Ճ�<��e �?��^��8;·9g�}�+ò��c�:	qu����}G������/{��1������vҗ�o��k�K_��ip��{�R���ruX������6�eYo��l"t��,��c��#��W �e�&ONم$��!�Φ>۹�.x
��U���;=�?Έ%&!s�>ܲ�x�"���:X,!]�I����@��.[�n\2
����;�`B����+��쿮QD�KZZ�A�A�A�Ρ�n���������;�k��χ�k�f����������@�C���n��G������w�VӵC'ʎT�sf>���}濧���F.[�U����/`�:���?��/�k}Y�����)�D���P�p�#�/�K�v⧿o��OOn"�)L=����F�!z�[x_�1#X���o�y���=��I�Z囦�i�q���+'1����jQv�8�
�!r�ތ�ʠ��)���Ssʮ̕;�d�5�`*�s.�����>!�!�a]yX�8�)g��s�H�w��L������_�B�v��י��-��.�9�����c�]D����?���8sϹف����Y2tAs�xг���`��lgi/ z"��ݸ��W�:E�hۂV�����Np;��Rt��Y��bT-�?��_�`R�/TvT���W΃&jhh0;�6y��>���h%8�BTS��''A���[����ql�kJ�Ā��P���%-�F��"fi��\N��7I?�U�آ-��Zf�.�7�I���Qr�L��#�:6N�y�)�F�eo�C��֓7�������4A��W�ͷS\����w]�_��|�%^��坭1r�2�m�%@Al��I'���h+'bé+R��f�����T�������@M�L�z	Rh����� �x�_n/�,�����R�
��2�vb p�(o���G�b+y����O�w�릟ցu�~�[��/�tE zkuDD��rm=�1k����LV�W�<���x:�hnJZ��Ta��b:�e����WY�
g�UM���`���p(^P-xP�������;g*���rzC�2�;ǳ�3'���Қ������x�:., X+��}�����O��D0*��g]�G6�	�ׯ�^W�fM�aV�IЄ^���m�Z�R
�D^�R{�o���t\26S��95(٨��\ɃP0)���� �eӄ�F�V�{�����o1I�g>j�0�}3
7�1[H�zI�� ͭ$�������J�*�h<���R��;U�"o ���~���=���	u����[��DU�Z�h��)`O��|�@BއK��J�;˟ �}�7}��8�M���N�[o�]�_�@��X���=��Q	�q�%@��Ҧj��,h@���S��]S�x���oR��Z$����(H߂7
�w.¹�Wm��a2�,5*�N��S1�V#���3�jcpvH����k�'�u�
��\Mv��,��y��25��/��ml�F�(�<6�}R (�`,�V���Q;o͝v�^C�v�'���*�jù��y�]*�GZ�`a�����!>�=�7	\�I>�ʿ��C���R۵��R;K���f��9c��F;��?�b���i�h=�w�3҈	�T\)NK��w�Hnb$(�����g�-���<����ȯ� 7i�ę��f�(1Mq�(�Y�ZՔH�o ^��2~�?#�ql���'yLaD�w��5 ���)�Ng�t�n\h��P�s��+�7qf&�_�>k��83ed-�fٱ�b���O�Nɷ��/���z��jۣ���lf�RFi���� =G6_����$����(��)�����A_*���h��B���偆�WX�"�V�/�'fcϞQ<
�,@�������Lj���\~/ioڗ$�����}�`���$.&���԰��B����n��/�M�`*�3��њx!ԃ]�j~�y$����X�T��^�#Iv#��.�ZE���9��
6�0�}Q/k��6��;`���pG��}~i�e���	�v�K�q�lwT���9����{N.Kpħ��?BRI-�z~�[=����/���w?�Ӧ��*K B��������܏��G�xS��Lc����A�eE�X�&9�,yZ��k2n��l=�i���l�� �؋Z�
jx���_6�Eo@��o�HQW(�(k���0�~/j����2+o-yB��`pӎeU�%���͜ho}TE�h��"q\���6�1>�:�K ��S^��Yt���9���� ��6$\շ��D	mg#��a�n�	 �p1 �;g&1�	L^�4+��ť�N׺��c<�f�w��O�9�9���[�D��noX��|٥A����:j��Mh#��U{�	u���.�^���茶� {R@�f	n��,���Q\��fu؍w^(���1�yѱP�s}�l`l��� ��چ��a�I��[�x�,�C|;B�:ȕz��.�jx��[lb�7�3g��l�����C��uH�1�z �)�R��<�Su�{������D6�B?Վ�ϭ��&�����W2�~ ɜ�Ӫ�C�"�=���=�����F�r��ɲ"+Mޫ���5��� 3���Z��Y?�� �̞��7/��c�4�`2��;��ЧZ��$|�hv�ϡ��N����6}'���\��w2�����s2�'�F�q��uTa ���M��V�g/��w-PU 煮�(D�:����è�l}r/̍]o�S���t���1Oԗjgu�� ڜ�u�˷�?�����7I.�Ա�/�������)�߸��Qaٌ^�����B��V�i�h�k�yf$f���6Lk�Ϙ����VG�V�� t��fc��ը�i�������X6Yz��( N�r4.��X��4�.��`���#j&����J�����$: ^���:�7�sZC�ޟ1�w5���H�x��VX�f�����.$O 1�(<�׷���R}]Yr�1���?�*�?����J�.��y��,�{�ư��l��3��qk��(�\Ň�D���^ܰ�����Y_ON�\W�-D��|��1�@��aB��bE�Y��k�}j�]�|��yK��J���x��T�8=�J�%�YS+��r�v�Ȃ3��U�B׫���l]_1w�}"I@9(�#��ߦ��i@���|��1y�[�81��贰kC�v�a7_njk�iWuš���؈'�`9��v�s<n���,֤���r߳����"�����E�V$M@�پuABw�0�e�xcA���!�KM�`5}b�:/���f)�u_~�=��y��3i LV88�w֘Z�X�-�]���.�sq.�=qa�����kI�l�"�4�{���Dv3��UC�WpC�!�z��ҏ�藀�.8�>l�1/��������x�I�2LΠ:��;��a�n�3H��A�@�����ޱ_
��;�,��X�.餜����ܳdO�?Ӕ��	Pd�,����s�������d Y铎��2���C3���A�sW����{J�]Vk����g?�������3Q;���U�0�c;.�ҠΝ9��)@�]Fr���H����-��7��{���w���Pq�����Y����]�~sMI)6U[�QI c��X�V�4:Ē5�;KXxd���� �~$N��-�y����(���h�D�� ���Z>�3�y���m�d���A���$��F�C��������vrE%/i�0�&R��XY�1q������'�v�s�Z=46x$(��������֊�S2n���a��ǲ����dt�h��+l�6X�'�����$z'/$;�H��U�Ȯn��	�QI��(��~�s!�<��]���z�nSX'�u��P��D(좓մ	M�}��
<h�s�M�|�M�-���������C�u��#��c ����B߻4��YS���\��������l��u)��1�m<��i{�SA�1/Z���8�f6g�-�r�͆��gj��ۚ��S������Â?��y6�����B_,��C�u�G���)���8��L~�'��
0,��L0����z���A&	p&����δe��V
lR4f�'�����N��T�qr��{��b�7LiQ_hbK�SV��bi^P�-dP��.۴�7@�z*g�8��9���+�!C[�����Mσ��̫���
�n/���lҨf�>O����ՒܭD�Zp{	Ó�n��Ų9~���5��Qs�h�q���q�m�\)h[�����Z�����Z=���nO!��Z�۾���f��`�D�Ă0%����fy�Vv�h��~R�l��2�����CHE�Eu;��"X��MU�s������ؽ�Ȇmnu&�^����i����ۜ��;qұ���pە�\%��[x���M�XhW��!D�k�7 ]R���h;����g�ߕ	<�R����	ę�1��2G����g��DA��o�����E��^ѕ����E.�vG� �P��}���>�-�J�SoB��>US۱�|�w��U��� ]O������%�ygԨ�y���y�[����$���D�Qt��c,1��B@Oe�+���Ho�[�̎�RXP#����)_�1'���|6��%l*����_^����*1Hц����V��X�n3ިk�{���%	�y�dÁw�0�玳��e����z%������>Ǆֵ
�,e�R�|2�x��?K<܇�N�5�'t����NLG58���ʿX �Rf�����"��B�Ь�����]Ϻ�{N��l��?���̳JP�U�`�9����"VG\��ve)�'͓�c�>]��c�����g>[۵�K~=�u��Y��h94ƒq��k9}�InO:�B��B'�չܷ�;�U��3���܆�s����%��U���el�g���R�0�4g=��:�z������4��4xCx�|9Z'���e�$v ɴ@�@B��6�'���X�f(��\ ��.�N�7rŊ�i_��z�[�=���rMFճ"S�G����n��G�ŕ&4�jT�+�O�U�k(,Ow_��������3(�"A���Z��y��Xe���Υ}��\�����_�N��߯וv 8�;����A� )dA�C��n�D$HR�t�4E]7f��>�x��QU4�oN�}���/�Q�
ߪ�˶-I�M^D��b��Xu-�8jb��Z��i3x�fh����_C��':41Mc'2����KZM0�_�VQ��m�z�%����SK��}���O��ˡ!0T)�"2E)S���p%�z6|w�LZ�T�n�Au���K޶'r�%h�d�ү'o�2�i��=�1�>.��v��aùd�m���f���S����>�����\�i	ʃ �@�a��T�k�.Û�B�^��¿�U�2 1k5֣�h�����z�@}��� F� �I֮���׻�u!L!��aK�Փ����~�![w�kk34�*�kn�9�2G.N�sIG7Ǎ�uM}i\������uU�caK�.$��/�x��ȃ��@��y�;����[��yDyF�K�ܶ<�9G$t�6��ƙ��GI�T�_u^�!�4��W@���w-z�]�H;8�exCa�5)�S17u�>�u!���3���T�B��<�������a,��ޠ��<�Kؿ�u��ۯ�,jͼa��b&3����{4JL�q&aSա�9��쵴>�� T`�w��~�_>��� u>��+^�ј|�hH�{.�S��*ww"p�D��m���;25
���C���[�x17�m$�[��b��i'R	���m��s�X�|�`�ɍA3��@Hhd���4� ^ĵ��No���C��oO��+on����q���x<2c�Cݭ�؛��ug�������Z����ƺ�� B��Jk���J�7̚�M�oFpO	��D��r���.q~[��ą���֕(��Ţ�B��`��F&U���{q�������Rl16�EQ!3�Bį����%�V1�V�L*��V�IpWN�xyHb�Ԧ�o��������p2�t�f�r�hT���f���ԣ�'�U���#U�5�Í)�?���~Z$-�O7x���i�h�\�Z@�-�(m��Y�+�f�uHK�����H������2�X+S��.=�q�E� �"Wb;����v������Go�g|tj^Z!�:=髞���/���g�Ľ�^q��̓�\����I����ξ�2%u\������t_��j������䩻y��\iz��Y�6�c�*�٬�Soj/Iz�Z�
\d_="^�������tP�����"^qizA5�ce�S�������d�+⠖�cÓv1�ejO0����O��`4���8::�����ÆX�l�|��&��zѵ��7K� );԰��_EEV'Dk�����3�X �r���zS''@�;�ŹFT��s�n��Mߣl6_J���B���_K�5�֣�Ԗ���AϿ����V�&oMy�9e<�Դ�֩���qi%Z��ǀ�$	�aU�!C�+F��� �XL!Έހr���B Y��YrC�������l��/�y�ڻ���_D�w�Hl؂���=<�,�^��b�yMm9˗=�䭶�3VSJL��uwB7���CpI��:#e�P��=�|gW����T�"-	K�V�1:7P�q��ܙ���W{�0k�3�60��U	���Δ��F�K�-���'�m�̨g� ���T.N=:�ig}��e�휹Q�-X����z	g�w��0�p��z9���Z��O��m���ƃJ����D�Ky;�>����=44�%z=���-�Y&&�찧�A �k\o��/ѩfGZ�R���/Hya�35�,��E�ڦ�L��+�2G	LoV����l��8��l��5��d����H�l
'�r�e�ZtL�mK@�~pf:�k7#�`�դ��:�M�U5�����&�̗����3�It�`\�E6��sF������f����fx���wws�_��<B�I	�uƌQ]�S�Jڅ/-�4Ui�F�J(�z�����0O$׉�P�_�Tvst���=}N��|d��xml��g�C9��5���!H��܅a�� ۷���y���Z��)$Z��VoTI:��M��1i�d�g��CU=ۓӗ�FR��cJU�������)�coR4{N�9z��R����Yt���h��Y�x۱%]��幜 ~�A�fʇ*�>��c�#zNoSaR۾r�nئ�������������⿲��ir�k�'��P�Еo��O6Z�!��穩r|��1A�5�ep�R{i{!'A� +ER��֝�"�����z7CD��j���k9���7�SR��$�TJ���g|���8��%�x��Ds��-�	^� ��Y��v���i�AH����6X��H�Qr7{l`)9��2/7X�6��L���a�8K�O9�J�(i�	���N��Upe��ŨZl�����������oqՍn��.�f/��78��zSk��\sv����J���gX�Q�Rᖕ�4d�À�M�Ѽ�N:�=&��^,���-���+��>�(y1�w�f���ҥ���G�ή���̙%�-3�yM��P��*đ|���pp�f'�w�.���!������Α��*��d�jހ���_-K�Z�&��p�{ߑ�ʂ��i�>k?١+���`��p}�TT�cq����?�u�n%N�l�w7*�F4M5�b�G�����&��b[!;�B�+���y�I�a���n�H�;i�>3��2��C�� �Kص��k�@�(�6h"P�5�Ya��T}5��3��?H���uN��T���W�ڂ�hu�����)�Ŏ-q�� Y�0,�Ԅgc������y�i�uR��u1�0P�Yy<������.�<���*3��G��=w,��d��n�V3�jZS� mZ�������x�h�^U�W<*��V#��l%=k1P�h���w���9��������o�-y���n�N�ru[������-���X�R����e��R�<�p�Ĺq+�v.{f��J2^�"��A��kC�;�ˮ�^��"�Vn�w���m���������/�ɱ~�8��������h�}�6p�����1+�m<��מv�k�{H��ڭ;`Vo�u (�YQ�R������wk�h���Uy.�s�&�W/w����-��G��~
_�ȹ-U١W���y���ο.�k/�Ϻv>�oS�ۉ�˞�dݛ����B��!�K�P{#6a,��&��a���(z�
?
���j�t�l}�%bl?�R�D}����L�;�׿�;tH����=�~q @�2z��$w[޴ROL���m����@�D�S��7�Ҳ�W�<4�'��C�\b!;�����^��2��L;�pܫ�8bA��`1�k[Ag4���IZ��䣒�ߡH*��^���}	�,CLe���mģ��^�{ǡ��p�l
{K�\X��C��݌ģ���5m�� ו�'�/�f�.dG2LUAu��۱n��xG����!����^IZ��nWB��|Q�L��G{nϕ�>�Og�-�8;�@�<��/����ieU���7��v�/�)0l�\tx����|l���4w��uf7�E�����k��QMK�t�5�ѵe�)���H��R;�0GY�����jo
c�R4�K��$u�jd�f�7%��'�L�u��P���� `�9��l12�r�|*���5�uB5�P��w[Xf��Q)��䊪m��fU��,s]�y˃�т
|�6s�8WV��<B���HXŒ]�m)��A���@�L��������d������\CJ�������A��XBݫ>v��)���.�Հ6rp=C�e!A���c�v��M�^ŦŒ̐C`�2�ߡ0���������ρ��h��sqf�:@#���o�E?9a��Y�>J�ᦍ+��E������ƚ�^R�I3�TO"����,��9XE*J���hk4*:�X�rp_��Z��J��YsQ�>��L�(J�u��B2������^��7b���K]�,Qcٵ?���$GK���K�ԫ��<34%��8�m�'�u~�,��0��s�[��2�J!b.��;_ͩ�d��ie��~����(V��@x;h�����L��.�4]��y̖s^���뾏	+�����0�`�B�|���B��~�?<���NF7�#M�@��%�X�=u�
��#�!��S�J�φp܄_��?A
.5:���ٖ�U�\��cruseM^UF��6�"����$ɬE��Ƕ ��ʁWގ�`��_y�ƞ���KL���-D]�C2:צ�y�*��/���ճ!�F���X�t��t0N��J+<�phLE^�I�-��"���
�>&��ֵ��7����:����=j�j�r��.�nx���Y�	�0�i�_�ٷ��K�-ʕ��ؔKe�Db�V7@\�n��a6gcSO���9�W[���.�<�(�)���p	-CX#�FS*$�d�1L�TJ�c�)_ 1���`��"l�n�&� ߪ�>�Ƚ�rh���M#&V�[b�	��qL��?�Qh�D���*vZ�X�RWd�z&����C�9�f�K�`n�s�nSz�匪J��E����T��Tᤄb��\C
�]7	���%k�%z�O	�NO׀6�6e�N���w�`Y�:J�G����2ra��z\�ynU�z���<Qc�|5!ٮ&/h1*�Kq)�`���?�fy��_pͧ��+�Gq8�~D�.]L�G��dI�m��uZ�bCsg(=����S�R/М��MH�U,�Rf �z8���9������ �$��B��c!��ҞUc�T0�2��\-(���y`�Q�m7X�t3�ig����ƑA���c@MW���)�7ճ+��Sy�$�.��e	qo�{5>	�8e��J@�'��âkn�b�ˋ�J�	_E�5�
��:טp�3��a.X�G/k*�.�B�D�Z�(LA���1'G���]9���I]y9��c�maW�K�3z�Q��/��O��W�����,K4wD-�h�=�L���A�i�	5���g�%&:)���.��)��l�k��D&J˒y�k�+t�ܢiR�_%�p��$V^6A�o.eq���k��
���+Ѱ�Q����r 
���K$,�T �'P_L��|�O���|��,8"�6$�(bT����qk�5��u��0���X/(,IhF�"��
m ��TE���xokU��Z�a�|JPaR#6����G
�	6A^x+ih0����KD(ϥD�X�xvӂN���x@��Lǀ=�@�\�p�n�K[���5ً�\�����X"i�r�:��A���L}���JS�j�����K�{�F��ݘ��]�����_ټ� �1�UTЁ+�����G*-]�����ß�KL�&����!����P<�J������6��P0�e\e-�|�#����I�J,�H�[8̩���A��;[�#�'���3B&�r�ս���o���(.%P�P
 4����׌3�\�ȸ�c�T��B�l(�ҊnX���[��~L��Ю�ZR'&����X�E`���3h�!�ZZ�Qc����ziBGǇ_֯[dj�ˋT:�R��=��YQ�"6�5��4��i�z6&%P*�)�*z,�}1ݫ�fC~� �/غL��pm�1���FT891m�1@��iY�7��a9!܌�J�>քc�$���݃��֜�,U�e��"U��=�φ&� =���T1Q�pQK���ӦD돏�����x~#l�6�����Q�l��d�LOSb�ML+��`�8*ڇx�w��2�o�n�e���ı����+�Cz��v���+�E��w��ΆҴ1�Ig_�����O]�j�n��M	�Њ�1�>�S�ĒOū)��)�Spս%�ԇG�1@�ɼ��"X�r��Z�y�sAx��/X�E6g�
��g�����q���P	$���5�ɗR�\E��1u�Xey׭j�R�`vb^i�ɗ�Ծ��y����s�m\��h:z��6B�(�+p<ؑ��O��]��ku�M'I�/��n�BpY��br�7]�bQ�ɳ�av!s�k������nq�̹%Ϭo!�Qr�qea(����B�ߙ�3�cP8��(�Ƕ%s8��.��t]/{3كXak�s�T�����aҟ���ުVF�ݤQw����c�񪄋}���¹��2>X8����޳�k��� ��	�Ӱ�;�������M�V<z�T�X���_Ɣ��WEM*���E�]�s7�<�E��g�qB�eTW]�=�ی�^z��*&�x���ˮ������6�ޔ۱q��|[���J1��[DgC�{V�(�����~lYv,D%~rGֳ
[x�)�_��l�s�FB8JZ�m�Qפ>p)~��/fF<%��R`�bI����Q�>�Hf�{���꽖��Q�Z���>���6)44��b�UK�dT���4��WtF��5Փ�e��S֮}�����	]QR�iB�X醟��VH�Q-��E~�N��5t[�f��
���ǣ�Z&�'ő��N��8�4���G��w�9��c�e^b\���Tл��.2�M��>4�n���ߩk���	PH��v���c�%�ۨ����i�cn��K��p����%2�����~��@P����C}�bq� Vl4\TO4#��:������KOmئB㳤t;
�<�n���vMg^��C(�r�_�,�����_=�.���BQ�Q˩l6����M��fd�X�5�
,7�N=�2H0���-[�����W^|�7&f�mޔ������irr(�������.��:y\����ܚ'Q��`�/�>����U0}�K^�`d�^���­֒��Hqǟ-Z^,��5��$�w����LR���sG�1��A�Qq�.Ҧy�|
rK�r�B�C_���0��P�7�r^�г�8�ԑ1�{���}��[ŷ������v���M��[(9WBW� k�oύ��o�,l�o�9G�7��&�S�pE#1T�ʒ�q9e�|����,џ2H�)����!��:�G���%���m���B��1����|�3�
��+M���d�if�)��A�e�Hٖ�Hp����*҇����6��hįN7����_�и�4Z��P<�f�E�� �`�OfU���M	�B�^��!p|Yv"��nv���&�5sN��z)�^L��l��B�)3�9j�~�x��q��)|�����̾�Dy�^���o�"�;t���qd��Ѳ��(.��-�Q堰��16�83����M_5k^�_gUsݲʾ��f�8A)�z��q8��2%���=�OK��	o�:�^��-��85q�:}��������l�ӂ\R���Y7�O�+���v ��b�Fиc�g�H9D3l(=���lW���ى�QA�˨��L*i����xĊ�K���LP6O!3N�������cv6���rZ�T�,�������A�\0A*uj3�����f�ce�LA',��8#�A��*��л~ߡ�n2o��W"o,ytY�_9�l{���T�<�Y��e�]����U�k����}��xa�Y��]9L[�]=���O��rɟ�\�<]?��eaM����˹o�@��(���A��^D�z�y�C��%��� %ē6�ٕ�?�Xe�ixk?;�k�xݟ�zLv�w���<=�VL�.l \q���֎e�U#R���@��(���$�L|�٢���Y�ټ�!����	z�
�hOɪ֕�f���Ϝ�0nM���pR�O\�Z��-�RIUj�O�:+�M���9۵)�����54R9���XRR��,?��Є���[kE}���V�-	�P�?�gc�i�4��{���`��p�C#%�\&������]�&o�t)䠻3�F&�g�����������CƧ�[5Z7J*vB����$q�Ϯ&1 �Fiua�	z��f���E@����8q��__b�0\�";t��[��I�M�G*�X����u����L�=42r��s���o�#:�'��M��_!z��c�>��׿'2���7�ᠿ�Y�O;@X���zQ|d�+w�qc�~ˈ�q�f�"�d��vX�Sq����j�d� vy��b,���fdr2���J{��6
��6�x�e��o���M�< ��SŨx�\w�%��~}�(G_�uuj×��������Jl���81?�Q2��Ļ����[M��zhY����jT��U���c�s��~���9�rp�߿$��4X ���ϡ$�
�?yMO`E����dϑ[f��=�Ѳ����6��^�����q{�����Q���QcZ\[�Aކ8��T"�)����\�Wt��N�W�Ĵ4;� ?Dt���"uy��=0�(��׻�pr|����m���4��OW�_L ��RQ �*���a�Z��yض�%c^�q�I�*�N)�����:Z)z�M)��.a�vw}���+ε�h@�N��B$�,�R�7xe%bJc�3�;���p��O��w�<�Ҩ���e2���䠣-�+d�U���U��.�BĢ\���|�N��ĉ9�X !�n����u��+Ue5���s�S}b��j���d�ك.��You�����̈́����<�3eA�����&�r����uT��R%�y��S�l1����؟l��]������V���g��Sꂸ�9g�^�M��	��t^9O�겫����ϧ׀k�y���&�>�Jbf����jں!���A�=��m������'AH��2�
���ƈ}�vT-�����:(g�i������1�ƻ�ѬΣ� $��T�s�~0�X�ƾ[�.��Y�9H�����A�cYH���tn�@U�����K�t.R$�5"���~��J�B��Ø��UY� �ߺ�h�74���͠a��n=�d��	��FOW�-֚��g:Qh����n��`o�G�=�.��H���`�1}�h ���z��7-9&0FTҮ��Љ�;����z��ސnVe&�`fA��a9�T!�-�y���F[�vd�4���,�yd����q�����wĈ�B�*  �=��[��n������k�x[ΚE�RA��d'm]�j�_��^�&1��,$H}O�+�y}]��p�1[+�N������P���αF���T1���ش@�c*��]�S�GteW��6-�o�fTJi�b:�F��+L�ؾ3熀��-��+��t�g�s�O���6�bp�H
r��t���&̕>Z0B�w3��z?}ao�r��Oy��#����^��7��Ǒ<����P�sl5d��n�&�齰��e �7��� �m�F����^Z�\������WHyL��%*Hڻ��"�9�����ϭn?�ߴ��Tx9� g ���E�n��D	�/�c�K;���p��3	9�c�׃�"$�:�R�}̟I��x���^�
zo�3��$��.��9Q�F��h����T\u��M���	�ߣ ���X����IE}~����W
��E�y>uM�^�C#�P��)h;��X�:`�Q��u�P�٪pv��Ǘ���Et����h������`k3�T��B3�J�雨V$�W���H�EI�Hј)h�����q��n
y��:
��<	D�����_x�]
P��t,+Q��:Y�xg(��(��h�q?���F�` -�Z�g`��QC�d��#���)�&��s�������7���ls*
KΘ�6�0�������fR�G��_���ڵ�Z����7���Ǉ�[@A<�y1k��T��;RJ)� �Sz��qAZ�^:����e�C��ٕv_?�'h{hJq��5�V�����W���D�ȓsjμg;֏��äp>eT;�,g�\�w�f��L�n��R@���n�E����J1��JKH�&h&1�\y��;܇S��5n�3�G�q&��F��i�������W@[���A:#"��G{r�X61 R���S�#gNKr������W��	�*�O�{��P-���=H������3,ǩX˟�=���u���,���zm5qX�2�J��;���[ݜEL�o�s�����:���Y�X�ޤRe���Q?�ܮ�5{m0�Q���Я�]�ݙ�-$&s���Bc�3��#�(I��i]3ϝL�gn�����_�����)�m��*��.�6���J���񌹙��U>��i<yOϷ><p�L�����"�����OM�[����d]!��m����6,�'�%�ݙ6�Q�[�D�'?�5Hu�L�!�?mߍ��^�'
׉Qf�ا��������i����|~Ңc�?����PW:	��#:(z�C8��9¶:���j`�Q�J1S�ř0a�/L�at�<x!|�T��9MZ�����1�*3��hy�aYZ��t? [���|G W�>q%e�q:+���ӽ�Մxۇ����x�|~�ha���,1�~O#��/�|J�ұ���蹾���M����1�N�R4��V��]�(�<���}��X����!��<x�[h����c�q	��Kl��F~���=��o�A����5��lB���e���E��5�ɡ�vJX'd��Q\yxs��jqv	[K�:Q�!+)Yw^9#�?g
���?Y��a�%[.$4��S�6�mkU�������Įꆉ�ė�Zb��t��Kֱk310���9�2���uLm�9^�ɖ�4�AkIP&��8��^��X�W�H� 8,B��ʊJ��@	)]�R�����8��(E�\�ة�,sA���➤Gz籝�}�6�u���|��WA}�
�L���b��w��j:�[��?e�ѳ����9}D ���`ɭ���Π�- ���M0�y�2���B��ͼ�x�5�f��폡
}q�����h흽�J2��V��&]�?�\��$:C���g��*����7�����Ą������"o���._�nй�O����O��ap�+5nТ�{ǁrhrUr���K�,���~ԕq5E���dȣ崩%��=����낝8J�Q���!$�=����_�~g�����E����-k@����ٗ��y�^[�01+O�6ᾯ"+en����n�4	�Y�^���	��ں
0q�Gig��[� C�Ϋ*"d�uvb-A�J����J�i�TĂ>��/^Dt"c}��i0�)���Zᘛ�s7?ڇ��mr _&�S�����z���r�*��(��r����؁�dܯA�.Mu~�1��W�1Q���"K��-�yX����.)i^�:���b�=��5� ��y_l�w�U1a��yT-FjBh��{�RbT��id<�x[���b�]9��!���.6ܑ;}%�F�j��VG(�\�������p�Jī̙tF!%��渚&� ��TQ�!1k�����,;Ng&Z�i�2a��|�J%b0?�Mx�y�|�z	3gM:��،�%���E�vaù�B.�[����M([$r
��=���@QG������������/�-���>d�?��su��✥;5�ֽ�A�,�O
S� ]��Wo`�[������;&�eQ���p�Ø���ncŶ���GM��79�*����]��Y�=������,L���|���zA��UB��rc'��?��]���E�P�O_8����Maj�	��N���@N ';ާ�m��,Itwgu��դ�3ף
�����@�'ܫ��Wf`�y`i\[�\1V��	V^���S���*��cB���6�5�����%'���<��Q�Y֪�P����c����[pks�]a�B8w?u�`a��t�(O>��Ê�[�}#�>��.3e[#v$A���tY�j��s� 	la޽G�1�Y�g	���gN�>M`z�;�7
%6��8�\q�V<
޷^r֏�e:���/6Xҳ���6s*L�2��#��<}!�M��ġF��� ��!��Mz�֭zHH�������Z���K�1豾��LW��C�Kd�#eu�����$/�;�qt͏S\)#��\�jJ�&b�*d������!�Ox9��"b��i��I��ܕ�U�=��k=���y/�~ut)^�������n�DLL���2��m���Fp�0M�p�
�i��U ��Jk�h �|]�&a��D1�w���PW��3���?F^܋C��1ՖZ=r޼��b�?�����`�	$�w�]�ww���,�C����݂���;ܵ�s�8����c쇽����YsV��}9|��@�g�X仡�h%L�8��)DPn�D��W�f^�ɳ	 MR�YZ�|����P�'��l���Cz�m3H3��7�19�T� �a��J�#$��5�Bd�����"e*���?w�0*q	?���2,��>���Y�	���P�MS���>Hr���R�n2lA�X7���7��:S��&=��&���?�u�~媍f!؊�l �>���n�'��H�Cv�l�;�!�� ]���7�¥�u��I$C�r��\�t~��{b�/!_�!�jϧ��M��F�4�;q���ʹ���������Oj�w���%_T t�IDi'&Q7 -E��b.�ް�s���#N��X6R@�j&������i��Y҆<�A��X��ٹ=]|hGxa�<v/��3$�!�q��o.b�%
"�2�ʌzR�D��}����G.���W��'����Ѱ����o�����c�!���F&�����������o�fX��;#?A�ߠ�7����kP��	H"���z�Z�1;,}��$i�����p5�a�g=���R"��{5�<�t��s+[�.Ǒ�)<����������9���o9�5g��o:G��V����ZԻGS�͛�,M�/�2���	��ق��Z��S����v�����潿��Y�ߊ�^*Z���������z#�BTouH�ps�� -B��[R0���&y������H�H��q����R�����EՅX�?�Z�j����Q$`�Z��Y��]���Z$âJ�]2d18
C-���Tk*�bX��LL�*)C��Fo��`w�Ucr�2�����]�5��D��2}���6�mxH�B�|�S�[e�#�KS����%W__�D�\���3���'&v�����I�᫲5�� ��Zܳ�t7VD|��%��I9��$d=�n�����s�96O`��嬿�E|J�ݜ?%�O�3�o�k�2���p�(gd|��t���W��0A��훬wKc)*g'y��),f��a��?��CC���FȈ4X~��"�<�,&X|����	5�9����Ha��E	Hl-lX�6�g���⻹sz��ڕ�X�"���=���H?��*d�3��;���ڜ�狒M��3�2v���J%ɲ�?�|�	�������k1�z�#7���qwE�ݠ�G�+� �r���y�ظ��ҋ�\^d�<��"Э�Wk��h��y�x�H��q��"���Bf�5�8�����uF5��[�>���ܟ���ZNP�}Z�C�M �,�0�2#ͱ�J��c�1|�[�o0O����I��o-��\_�j-�wMt���u���uʊlm�WY�Nۺ�#D	O��2Z��8�T���}����!�盥n�o1����>���AS)\���쟊Ԅ�i��l��-]¡��M������0,��2�w���(��
���OI�9@��8�/BZy�k���g�6��AY���Qes�!B���ؕ��~j7Z���F�Z�u�&�E1��n�kJ�\�D(J��	!��i�I����^ܟ�_��{�T��dR���˟���"vj�J�S&��.c�Ŷk�r\d����\nQ�^c��w��IAi#Q� �n�=?U�@�p�o�Y���ƅ!:ؚp�������X�6�v6Hd�#�[����ٔ��0����`��5L��F$�T�d�0�·�h`��M�Zޣ���&_�;w��er�����UZ}���I�s��B�I���2|��OI(�f�M��Sǯ�h}3X��A��j�O�K�N>�Ty�_%�������"0��9�٦�H�����dl���f���@�#o��Wd��{�^��Ɣ�]������;�L�	�M^�Ǩ�D/B��!���)�~���@�?>Wݥ�]��)��+x*��eڋP��>^8��lq���[��&�oS���c�V!�1#�K��8[�E)��t�-;6�'S�EC��RWn������ޙ�Ɖ�#	�kof�u�x�n����=�l͒�^y�B�if�L��wE7_�reՠX'�3���]�7jqX�<��F�c� ������t�{4._�����/k���BDǌW�QQ��+��gm�ōW��������җ�l�yo����~ͺ�^@���T���}:�;���k�h<*Ɗ8B7������~ʫ}qo����Ǣ~���%�z�Ka�;do��T=�!%O�c��#����<����;A��������vU�X��ޭ�xqu�r+> ഭ���lw [ԝ{q>S�?���k+�?Xy�{����7J�	�ń�
T�!]�d�-M���Z1ז���@5�Ւ�9>w+M�� �	w6�f�?��:��^�	��F�6���b���;,����_;����	���N�P��s��E�od!�/ڦ;)����MP��l�9kqK�D��e�t�4;�.�B8�JX�a�~����~\S��5�7�ƥb=@��V��s6۽u��Ü��w��wWO�s���^�	5��%$n�(�A-��bz�h�D� /��g�l�U��'��*���M.)�'"���H��x;/v�Ȑ&�^�v�7�s���I6G��BC5~uf�N��e{�K1^�dܛ�<���13<>Ta�p�	�D
MU��`����0�d�{�,�b������V��y8����?����57���m�`�_�{����ɋ�ԫU
��,��ު5<����A�0�]�I���g8�	�f#��IR��%gyj��������a֝�>��Eޜ�j��Y�6��v�z�|�; N��%B�Af��A�oS��ԇE�s,߆Z U��4� �ݽ3���E�_�T��]�\�?Bbk�:�O�clXR�N�=��*D:�Y�c��t�B�s����tpxx>�_Ͱ����U��/�4whoew���G�6�X }���:AdP.G<���������y�T⏲�a�����Tz3������W-�p��h��´+�}����[�K����n���hj���KO/�5T~YX�^[�٬�Z��	C�ټ�e�}�h���hv�cr/����?
\��� rc���6����+K�����	���P����8F�˚��*A�:ڝ���ǩ+v!4��角q��d�'^��h��˯ƚF��k{&�JK��Ad���,|���p���Ij�۠�z4��Oc�[���9�-�#�.�"�? rIH�es=;�$���IcP��$��bWx{��fٵ�P����g��,櫨�������"-������o�=�Sܝ��*䭕q��(�{��2	�}!z(ZMz����o��V�yu�٤�jD��|�H~�S��ʗ�C:#o�{Y�}9I�P�d˛�� �Ǐ�BP���lY�!GC@!�'��t��e��:�� r��g��}[-��zZa�g�~�d I e���07�Ak�1���$�I�W�EM]���b~�t8۲�"fIB�0�
(�s�un(ם[�s�pZլ���٩�Ƨߧ�}TJ�����c]8�cY�_��h��gc��,���:$nK`��\%cd�3^S?�\xJ��ZCo;��6��K�����q��D#7QW���sP�V�f��|�p��>j���?({��|�AG��؟Z%T�J��8�%e/�:H\j�|ը�Q���5'�9��L}������(��~V�cZ���y9>��o�[V�W�Fw�h�[���Sܵy�?r�3M��&�.H���gN2 �,��w�t����E>�p[�~�P����ŕ}������5`Y���w5}@��\���!�۰���]^�0*T&�3ê� ���g�<u����p�_�Ly�
m$Q��s�
1G8��x����`�z� ��s��/|�^�kI�(�������Ӷ�Zhk߀�f��+����p��F!�+�|�]���
��]"�:�+d8���jE���Z�x��l�Uw���>��E�M�h����>��A5,[� !m4q�i^֓��J�1tYV}���X����L�fpq$[!����@$S�d�P�L��?�5-yy+	E�rB;�"��͐'����>p�w�5r^��F3�i�^&�U�M���?�i����6I�r ��%i�mo�a�^P��Jl�";�s��F-.Ր��ɯa��%�/��X=#��MX����W20K �Y�`���=�b�>צG�t�m���,�5����v疜l��]���I��r%�}ｖ������	� %�V!����x�a�9a( �}u���Y_Eue�X?�r�h�o�x��W�7U�j p�boS�v>�>5�z)qt�YQ�z��:����wXi��h�[z�`��ݝlhB��-���K�����-�G�L�_��wfn3�/�20@L�hq�X5^���}�]h��_���N�@b�P���wCFx n���v�{$G�c�*�f�����*���i j�����Yw�gs�*յ�ӵ1+���D�Ւ�g����q�E6z3���T�!��l��������`��$�$��`�&�o��OK�p���Z���%@�Q���A?�tY�uU�О�u
�����@>�����l���`�Y!�yQ۞˽��KRV�X��������!G�2�N�B��I,z��������vp���>�wh�|@��Iq�ic6q�8�TLZ�8�G]$��슼�'P:�b���ܵE[�Ƚ�x�r|@:���ޖ�C��!+Wj�eHZχ���Ψ)nB�ic>� ��Zimtʝ��		�t�V9I"+<ʿI��(F��%`�4 W�y�iP��Q?�	��62�7��iϽ�������AG�"�R��Y�@�gI�Ԑ~>�=� �빾����*��?C�kk-5p�_��3!G�ΐ|<�#�_�LA%mS޼��������>$isM�V��oWzْ���.�<!��V�B�sʌl�b��S�/Ͳ%[r%�B� v9A����:�B�B�fh<H��T�y偟���bF���NbE�+C4�v�Ϋ���G4��|�2�':0�߿�"��g�Y�ʇF3��ص�T�~/�@wq������$���2��:Ǻ�6�v�H`W��C	P�F�
�xs^��0���� �5�Q-��D�ƚ���}�ǵT��!O��&�y9�������[�pmbQ����#x���I��mbH��P��	���Ω�rd�� mj����μB������-y�F��[J�F�h�u��M�h��N�]���t���'k��a����Ƞ�S�đ]�*�ȑ�.=�w�L��$�<�*�Z8�H�]W+�qX�0�,�l�3�.?�����O����xu���²B�{��"ܭ���JW/h���.اi�QH�ѭW��v���u=8��:��
4�ï�4</=��t����Wm�.��V�7`v�c�Zj���5�x&��4�xM�B�-�����*�����p'5����v�����?�Û�U_��;�vc����Z�ݘP���ϋp��6ߋfux���-�S�	F<唝X����}�h8����Ou�K4,�V^_Z���
	���葱�������y���<�L'����`.g�uz��>Q�o{�ؾ�%���\ys�?�(ʭ�?��Z[yV�We�ma��~@:�ii���
S�|�+���<�4 ������I�m�7�o��Q��N6���S�Z;$7�����H&L)p�\m�i�q�����3�f3�� d6q IY��ǧW��3ش8�`�07�����=�j�ϐ<p32�����}�Kf^t��#�3,|R<�5��F7�a�yp�QHKR��"�"JT�z<�b�Kպ៷Kr���]�m<�Un�}�Z�gis�B��@�)p��)�.��I�>R����'��F��-F��/p&���k5��*%E�C��}�=S�u��e���Ix��"ͼ7�.=�N{.s^�)�t��ng��˩m��	�9�(�?��Y#������D�ޓ j�#�@f�R��;�������
<{uד�y1_w�w��P�j���U��>3��R�)���	��co��m�,��Gm�����Y�i�KW�f��p���$�� t��U�rÿ�MZ��\ң �ɐCX��	��?3���?�B����kPV�b�n�0d�+ �J��6
^6L^2�����Y4'�4�é�x4tY��|,\�~�M�a�2�׈}��|)[�oR�ȟژ�혠�Jtߒ��kWu23�	�Mnj~��֑� ��݅�j�eF�Bא�ocs	0�Z0����� ؏MM�](�� oŮ-S���|Y9���<�������z0�_����V�?���NCag�"L����ʼN"��w���0{tbƫ�b������w�f�?pϛ+
��bãS0e����'�adS��rm�
ŭ=�G �B"7�Q�^mka���B�"��b`&+�)�K��?�Q�W>�^w�2�u�mĳ8RR[⎨��^����!'$�3�>/�[]�F�9��y�=Z�L0C��A���l�a�i���N#�Ɓ�Li�d�⫫�/.S������a/����HO{H���Vq��r�P~��ⷻ;Ĝ���z�k�?Q�McИ̩ȭ�3����-�cH"1W�?[�4*"���Щ�t���۾OM��>�Z�P+Y)�K���Rt�R��X_����q��[zpr;������O�$�OCe�ͳ��+���e���Lv�W�B&��Y
�+\���=�|ǽ~(�<�^�h�A2rxé��;߆��m^�����-�jܜD(�+2��ӠE_s�ũ���{1�m���P�����=ZN��"`�mY��a`��]ǐ��a3�����ov]S�V��1£��w��v��h����j�!a8kr�Wa��`a歨|՜®*��[[�2�|�HAIG�O�N� �D���'���]�YY(P�1 oN��؞*N��mP{�.���Uy����C3��� ��U3_}7"����-J������n�>,��`D񍉻��f|�G9O�<�I��vf��	.�̷� �I[|)W���z��o�w��5�\Sw��9�R��S���D8�D"�'oѵ�a���LR��xi�Z���0H!Q��9˖�����T�;���E9���&�~-��W�]�C 56�]�tn��oz��S% ot���*RԀ�� Q�$9��;w�	!�d�3_��f��}��I�⌀��:+�� {F��d�i�;�� �����_��7U`]X���%ے�9
j	�P(W0�`��z#M�̮}���Q��L�l��7���L�s�=�7�e�G�o�
0|���H�Nv��f�4��~$h�-��n�z��W�Jo֬�Ĥ�X�l:�Sɇ������<O:���*���]o�S�f���g��НT�t�����| �X��5P�
c��,�L�ꅍ�J;�mZVqjE	�3�ē�ܾ�R�`�9�2F'�Ze�]�;!w��ㆷwޕY� ,ɐZ-�|uR�֤���U��
Y�ՄC�,A2V8#o��8��՘]��y�z��d%ǋ�0��W?ڿ�ا����9���D����l5�vA��-��L$��
ϴ��^��/S�\� I#.�# b%����=v����{H.h��c]�Ez�GL��*��3$�h<r�����T�.�>��l(��2���k�Z� Z�����v�p"BZ���,W��p$a��
i�Mv����2~���t��9(w޶��[9�^O[0sm͵>�QW�.p�y^�A�w�����O���7U���h��ߊc+�F�<X��|�=��E�B��S��?S�V�8�@wa�}�X:6g�Y��|S�0$���1�"HҊ"��j�z����Y㬫������{�fL���dF�4��"a�sSV�Κl�ciץ��J�Lyv�պ[g�D��I��Я�p�p ���Qɀp�˄�]�G��4h�Ia1u1�>;��%���n6�
.fW���J��<oMe?�TC�9�5�:	�I��<?��0CJ�2	�E�ZÔÚ��?#.g��]��eu�q�x���g�����筻��&�vͥ��q�mV/���`� �S�ۄ\����|��E��l��haʙ0�����/`N�	�T�?��Z���1��Lg]��,�6��z�"u���5f�
�Q@�z(�I�z�5Un�T��`z����&Wc9���|$8�:s�Ń`��$y�}����0kn������'� m}����l����D-EH��b5,����_�6���eGD� N�T��$�F�=�iS�z�
P����hyr�}�)^3�ʪ�r�c�)Bai����R^�n.ykZ�2�rD�>ѩ�cAu����W�q�7��m*�����M���s߶K�yn�J�GL��=r�g4ZW��r'�� �fnH3\��s&�׆���T����%���Y�~s��(:e�媔@T���qA�Ra�!o��fZ\k@aƤ�f�Gd���r)DF�;�:Ëo�8o9��t�b��=�о�p�ĶQ�R��v�>��N3ҹ���*�좖P�g�
p��O���;ۧ��y�I��W	jӛ�-=\�t�h�l)P]7��w��~��0ԁNP���¾;��{�����j�ƪ�������R*�ӎ�t�o�R���lL�?է���4m���k�뚤-�R~i�7�$��Ӵ����g8h={�N?ܑhܴ��sIH���V��M�V
�+���{JC�sBfst�����(2 ���gj��LՖ��۵�+k>�G�����T�ʗ��5@j�מ�h=г��f��A�K�y`>'���Iǖ�mg":E5qf�j��z�E�0���*�s�V��.p¬���=���Ki`j�,9y��FCan澩��Q#U�J۝_%�<w֯�����P�iz��D�0��^�A��	5�� �2p������ϰ7ڵ���gM�Uz�d��O�ل�R.@�C3�kr�N��"&*:S����8��6q"����Փ�R�`� ��Y-,��v cU�}��K�y��k�E�A��_��XzgN1��K-��]���Ұ�:��<���g�߾X�K�v���B�T,��r�<oPZn8����hb�do���O�sG0^A�_�Z���z��ӞҒgiY�Eߝ�����m����ފaI�/`��c�ƽ�.P|0�K��+btؠ�Nu]�L7�q@E���3�3�ψ�J�;6=�a�д|U�dcǚ�z�&Ua�)�q�<+���̠��mc�pZ
���P:�H���.}�Su�wHk����	ޮ�y/��2<uMGUG��x)[lHm�(��o�e����M��>���D��G�jC�o�Ƶ0*�A��_��2�PI���)kf�3)NG-\��N���v�)���Y��������y�[[;����i�G_}=�,�����*�����ۣ�Au��De����h�Һ��)\��k�CB�]��'):㏳Uo�ı��3K��Z_�8��-I���m��8�y���n5�T	^�D�����J:1ia�j��q�K�ʡ�˹P��F�W!5�ƚ����4�{݂u�`�y��f�OPe	P�+Am�w���a����R�T�vEZ��:2���)��b�Eճ�G:+&ʭ�E '�}g��%e���灁�R+0���Fr�~7]|q-}����s�y�t��r�U&�:�?od��/���.H��'�w>@@��jb{q���f�R��(�-��?[V)A���s
͒�m#$��ri�Qk4�}~�M�ӡ8YｊC�����t��;ȩ�g%�q�ߡ�K�e��N\��A�7c���?�R����Yv�j��z�)����Qj������n+�d�`�2�7<9�O�����+�kx�-_��tŗ4h:�����7�����徣k�\� ����0d7H�*��2��@����;<* �1	�?��:w?���|�\���u�]�z޳�u5�&�/k��A�ɬ0'X'��o�w��v.��PV*��H!��)��K��j>� y$B��'9���XRi�_G��Æ�9��{������t8-5��N7ዏ��C�����)�6y�8�/�$V����tpJ3���_��:�9g�����A��h��?:��R[�O�8]U��톳��$9��^�E����bR1��+g�ݜ���|Y�m�����R���M��ŉ�ʘR�R�7^pR���U�A�tzj����L>��3��T2f�LP}��}�j,�r�~b�|�o�{��&���?��UO�j�ڢ�)��z|�%+-�i�UTSR���3lI�{|��#�X�D��n9B����PYWY�����@L/o�����)-�S�H.��g�yg���W���zl㈌�i���,��%�6��pH n/ܤ�w,{P�I�m|X�uCbּJ��2���.lA��wD��ձ���}_T�-���A���:tt��S4��&m[uV֧�Nu���A�M�"q��g�����l;h2UH�ˇaY��BeU�IƔP�?y�I?�Ń�3[��{�q�S
�����~������4LA��8��z�#��N�+V
�����n:j1.M����%ʀV�*�e��Ƈ��J�k���^>�}�H1Z�S�%��oBX�d���a�{�U8�^3���#�&�A^��؛�N��/�,a�ј8w|0>(�/5bQ|���WKB�U(L�C���ɜB+H� <\FYbݵr����;�U_����[�R�7I�6o�M�����BJ��m�U��'�9�/��X��kb�+�5T�E5��(<�~p��	+�}�Dn"�[���b�N�zc�ΊYv�ڙɛI�,��[���IH�Y�����̢�y�����ޔ��g��*O	�'��z�_뷭$�rJ��)l�	�֔�	&�Zh��js�T���Z<J��أ�D6)�}X7K֣F����מ;��3ũ�-V��4h��o�5slɕ��1�{1�be�"�Ңѷ^t{�t�Z�V�S��X1����Y�m���PY��@]�Ò�yR�q|4�E*���#�MQ�?6�>�F�n�%n����_�n��'] o0��H�8����A ��ؽ�\ˍi4�!>9��ː��BV���G6[$S��Ä3��_�X��n��G�O�Zڗ���B���|!�'C5y�irk@�S)7umУш�u^�>��`YO�A]�"��8�QU�0m�x�}��LTǌ��/�c�-���s����D�81�͗��Y]����gC����Ӡ�D��M�}䓀��S*�Q	��o���̍�Fb|�D�|n����j�a��ϼ�@�^9(_��CQs���OM�o4��Z83�"�E������Gf���lN�,<�C�`���e=G[��L�w�?̕�˅���m2���C���{Վ
��h߮�2=�2�BM��8���cR��lz�� z��f`�ŀ�Ñ��wB����)֡Kq�gL�l��"���U�Ht�������{��:h�|UW������a���=]]TJdg�M�W�j�,\U��ypk�v�}�����M0a�2�'&�� ����%Z�-"IOQc��`� y;���\�>R �-�T��*
��-1��޻��F����T�tx��*Wz��v���t��a~�l7߷U�[���q�O-v&&-.6���X�nY�Sɥ|��R��:���l�N�j?t�ɥ5�'vm4χ���A� /:[�I�9�=��
�/s��O/��DL]c&����KA-i���f�y�bn�{�UR��r�ڙ�%�C>KJ�Y�K�=��z��\�褥�}J�����a�e����ѡv��m-���c �+{��A�ɱ8Q���^S:\z�hz�_g4zё��x�aH���a*�L?���M�c���.y*��7'>N}FP�_C-����Qҹ�W�^�^0�ND�݌>�@���i�F��W�O ��x�$H�f��~���>�G5�H?{ �C�S(%G������٤n�}a���M�����@ӵȯzs����eŭQFFP�~\�;�( X�P!�
d�h_����vd�җrvx��`�	��X���[���GZTK�����UD��.�~��bA��١��Fx��j��@�:�L%��c�����gX�d��MT����I�Mx�!�S�bc��:��x��/&%�z�R��ǜ~���8��.�}0��3�*��Q]Q����롕�i�?(�͞x��p��.�6M�7����i��A���Ov'�[�ࠟ�n���4�56���+�AP=}�c�F�6��כ�"��O`��e1ZKlt_c&��?t�=v��D_mh�FA�Y�U��]�H=7�'�&$���Z*T�w������� �<�H/�IXz�"�15�g͏�%B?�U
��(MܴGaZ�NNP6���+zzY*��[x���nm�<�_G����kt�����*B��o}Rˀ<Q�R�3�m@���$�/���3U����U��p##4������������lMD�$�sX�gS�փ�Ź�]��A�z�+toK7�e&{�����]�~F�d�0��Ι�c\9v�KH+���gU�U��o$�Loa�����4t��1]ϼ(���(�=_��ٺpOHZP0͐���@��A�;H���,��9PR����k��q*D�r3T=��1�k��k�i7?<��ۯ%`� N;�,S%�Ł�Y�ܬ�i�r���bG�A�mCL3���BD�|�<�q`#�W���V>fd懸#���#{J�5�0�s��Kz�Z6�j��s�N"���j�//7�_
���So͓��&��[�b
T"	�^&�"�7IB�Y~���l�\
�O�q=#�����I���O	{�_��I�k�A�ȩ9�b5ĩF$΅���e)s^A���лT���,�h� TdF��*gn�pG�<���;���1[��W�@~Wԝ�^�P�^��D�\ș�%�[���<���փ�̂%\j�J��jk+��q,]'5�#�C%O��a7W�̽���|'��e�y����91�y5��s���~��m���L�RQ F����W���E�����'�S*׳Җ��@��Y6���r�v���?3�V��&���[��JI��P�p����Ђ$׻���]b��қ��F�����y]����l���������T`z����
����#�q�O��<��z��-����t�Ɠ� �
��3j͋)APW�4�'v�ѷ��F�1��mV����EN�)��@���ǟ*�C��h��c�����f�3��[�"�����耠�z�Ԛe�	�>U{9 �@����R�]$��	�xN���rvk%��]�6�U���p<R�^M�Cի�&��O	��S,!nz�T�N��ɴx2eȋ�Z�0�w�����%�)P4�<&���&��=�|R��Z�Lc�9�Ϫ��f��-�p#�/�����< ͱ⚋���0�!��Ixo��H�5�T��K�v���O#������|P��=?���?��o�-Y��4V���LǕ�N"�H�V '?yN��[�������Œ��D6=D_|]o�,�I!�v�`�8���
#��R)��Q���dx��g	��'��c��˷�]x��r���x���A�*�q�OjZK?��c�_�C���H=&\���@�n���}5�H��]_�3|�����-�"�~���*�����[�'�V�b�j�o8�������b,@�6�V(���:����Ei[��հQ`쩥+����Fo��v���jD=��(�$r��S��އ\��⥈�rH���̈́sz���\�1���8@���3+���U�6��B4���� ��t�r�d<����Fw�i���G��#r�/�wN�JXriDH�~�$-���w4�	h8;0�b�c�"$Խ�d�T�=�?!�Y� 2�y�k�� G��%�G��(3	/��UzGvwH��f�s���]��p��G�j g������{��
qi6t�����#qkS^��2q� VQ26P����v����ٴ����~�F���j�7����TLH���Sf��ZDC�1����ag�M���}ǲ�:X��{XAe.I�� �Oz�
0L�G�X)[���6Ǖ��,������G�&��b�*]=�t@w.I�dB!bo]������L�q�mPf
��w(qʼ�?�˪�|P~�)�d�?�Tg�2��j�	+� �	|�з�Q���B�$%�����)�b�Z�����\���R������"�b��;�c�J��	�:L}-F��ܦ�3���21g3�x�2G�6-��Kе�W���zԎ���0����Uszq^.�͛k��8��:��k
��>@��w����Q�q��3���YF�JV���^�r�$�W��9��w�6�pf�����o�E��G�;��R*�9�Id�3�ɛ,�%����A��a6c.�0�ς/��Z�c"?�1p��1���Q1����X��9�J�_xh�h��̏�c�0� �*`s�iE�V�&�5�0M�?0���L �9��t�ݽMn8,-�����=.�/�W���AM�F����Lg��Ct���\2s(D��n�t��|��-�BA$�ٗ��;�1�I���*F�a���uP3ɞՊ�>�R���{�����0��Q<��v\���g�T�֐mK���?p�V�e5��6�і�B�(�i�H�ٗ�V���}qLs���8�,���d��R����	�c�Qj���K��5����h�g��S��"��{v��_gf�P��F�$���~��yw��U�X����:�_SO�݂��Bm��Y�$��˄n�V�m� ���7��}�P��S�sA��gL����K�sˢ�zh�|T�:(#�go"����~*��HN��F��q���!;�V���y�f����(�fIr�Ɵ���vq����.a�4[�y��[���Co�A��HԧIu�}2x�|�$\�oj�O�UZ2*`����
xH}0?"
k�� 1YuK���0K�,f����kz�12`��������[WF|��O�����q�Q���V������^�a~��滞����[��y�/o��-���=���*OM��2��^~�V(�R�07`+-���w������j�N����z�+HB֞zP�����`�m�r���$x~�����Od�au+�khR����n�6��Z�̞����҄(�n�]��%��%������">����^aϊ�u��kL;G�oP�Tj�0lf�E���I��SVS_}T+d3A��j@��̀�l��8���GL�Hi�ƥ���\ƕ�����O��1�����;z`�!
Ƨ�DP8}�*��)��XӴ��fV��m��m|�䫗=w��C��a/4�!�v��gذ~ߎd�j%$X�x��}Cuz���]��Ȃ�/���<2��]����Tz�rfa�L�ޫ�����a;�'<�-"3�n/&tǂ�O��ؿ���ڰ|�lGZ�AH��J&�#�8�_�@�,��t�G �����9]����,$�����C�B�����E�����i�{A��;a������[��%K�+1�����̾����G�t�9zt��v� ��p�+Q�X%b"����gք����%����d�|U��������N�}Aaa�	K����T�V�61'�Η�N�z^U�$�Tb�[�^���:��f;�����Mߺ6s�+���sVx%����R~��j��'�45�Ld�B��w��o�$hyq%^}+��>�-���<X�L�@j7BG�����B�&�W1�ä�`6c���/|����p��0��!0��v^�&�2d؊QOQ>�.��ISտ��`���H�NN*,eO�+L�q3�+��(dW_C�
�|���.:�S�p^w�֔(]��s���̖~}�J{�����;1���SMA&��+;�o���q ���)���)�Jk�B�
��+��v���]�N�34�|q�� �Ȏ���V��:*3�ˇ�I�/�ǹ��H7�O�����|G��赜��P�v8��:k�b����FfW���JR �v"����q��V���ò|��R	k�(󈨤�|�a��8�
mB��vgR��ł����ι+�?��/�ܸs�"��]��,]!-��7uY+�K�.TN^�l� v��	�6(��������p��d��3S�9��1��	O(���҆u�������,@U9�P�X~�=�S=E��K�}1�%g$�{��V9n���n�TE���/�~�P�ג�p�Hf(���Ug(c���u��*�zQ�\�Kt�{zf���r���&�Bx�y9SL&w�y���61{5��v�-I��E����i�hV�)ܶ�~�. <n^������W��c�ܐ��BHW�r��� ����,�;wq�
��,���xם,�:����u��T�[`06M����U�ůEV�)�``�KΉ��XU�ͱ�����p�]+]F���>/:�}i��sLZ���6CJP��!}��k�̥�� f��Z_�Ӭ�M��Z��JʙB��#[&���T7>(d�4��Eyl4.��죦a�R��;w���Q��ZŁΌ�yX��Ņ�S���Sj���`����i�ȶ�>���dz+�ǲ��gv��=ߊvf�=�I�-oM[�G�#�;+�t����U;M_���%�Y8�/}�[;CB�6d��݌?��-��Ŕ��x����5�zI8`,�,1�q�4����L�ؓ'${��V����w�N���x L�ևNw��Gԃ�c�3��U��B�OTOĒҢ~��aIg����e�V�cB��hUEUz/�.yB�ٻh+����0�l6�,��}�޺��T땹���fIY�A�����2�2����͉Έ��6�c�(�-�r4�X����.:��R����a�-����naH�%����-�w����!wi�qk�����~>��xO�z>Q��5/c\�`�p�;V�窌=���-n��i���Z�3�Qn�M�Pܒu�Zo�t|�8��'��M&��}G6J�̐��/�����x��^4��g~�������)�	��v'b���93Ys��.�+ ����	�NϢ�t��x���W+#�cܳU���+�� ��G(,�/�����SM�wr�6	����M+FL_��w��[^ÿ�U�ٚs�>ʸ��
����6��=G2p�uՠ~i��FΈW�b�*�0�\���:GV�*6RI�n9*�v/T�b���b�S�!v���k�87^p�a����`���Hk���	���$l���Zcԣ�į�4|(%�`�&�܁Gڌ�qŜ_�Qt��K?�ߩ惡Bm7�u� �R��3zޒq~Y���Ϝ����L��I��'���^��k��`k�c���k!���>Ҩm��l��U�o�1��iU���O���C�BV���ӝ��T��n8����p��Y�*�Ӛ���ZT�-��y0?��6�\��V�	� ���@��BFu!�/����'
Uv�%����q�K��t��W��]F&���ȉ���n9�]PG��J�U�Ȫ=��޿�3���$@>9���=�!x��pW~��V����oYzoa��`��r���C�Gp4�UR,�8du�.7b⼙��C�������a����&����w@���5n��ҡ��_Q��bF�j�Z]��H\}��aB�U���n�!�I$D		mo�?ӯ7}|R�߃?�	C�/�׳�x�����jU�ցָ����Co<ێ��oړ���J`kߔ�0���-�VG�b5�+T�5���K��r�{t�;�S}wU�hJ������-w�O��r�,�u��6��[�������o�z���D�2��vdQ锅�G4����Ʋmb�_�S'�9����@�@y�`�i���$~׏[{G�lKJB��E��D���EK��6P|�^�r�v߯�f��c�q3M��Q��!�U)!����Z��H��GA��G(�.�&CO{nd��-]��~��eK"�����)@9ߢ�b��F`�Æ����سS��;��*S鈓B|��Wce�!��/�|�\�,��kz�w�B�:k|0Mt@��AℏEu��K	 �8^���E��.��| ��KՆ�չ(ћs�˓#��v�\N���w�u�<�l�_ψ���cj�bV�#���Va��]-��Y����F��ّ��\ww�D��x����8�=���M?v�@����T����OV�� �������$Q<r�[:�JU�\4q�[��e�68�~���4!����M��|E��F/��-�=-���X"k�ϒs��ޭ��+��?v"�\��8�����s%��<#��`RZ�Kΐ� [J�Z�U��`�����L=]�ss�?�fpo�����㣌�Z��bp4Eh��BڜEp�4R�LG����{~�0J���m/��_��X�cğ\P��M>#[m�iE�O�}���K>W�w\8���J�g���!���}����Q��q)�����E�5�E͢�µ��u5W��CD���/ױ�zjt]ӈ�8�bF?���׸sX$ e���.)�)kF���MV���H�d���dI��'A�^�P�9q�z�'��topp�mM1�yg�p7��.���U�Ǥ���9t�.F�	U���5Ⱦ`A �	�a6wk��50��vw���V��(��Z�!���&㿦�W�]`y��q`x�iγ���zz�\^�(���S���[�5�T��dC�ײ$i�|���nk�߳�%ϧ ��;˝�ErY*��Ü�-��
\`�f�x���l$٩>�@-u��`�V��E֑�F=�)8��W�V����c�����@�!6�����A!�fk�p�2�����or���6G��L�����\%f�k���/�>� n&y�+���,�&Q���պig���`�t� �͚�t��zE�ᑖiN�>Ć�M� �]�6�C,R7�9ݣ��l�>ޫݒ!��Ea�W�0�v�*�Ҋ@�6����$�:K�&�� 5��� ���DB�Vk�;
��	V�+�p��	5�R[��A���7�z	� xˎm.�e�L�a<�% B�Z>���~��̔t�(��MC����X���q��^�gm1Dr>=LCϪ����-��i"�f�S�9sC��\4+�ӻ[����P�SQ����7�Ï�R�di����&�KY���[��\���ٓ]q����}��J*��qI��.��0�F^��u���pmΦ��������>O�qwn��qq�1��U?�1�P[�+��a,�.	�v�Ċe�?�~����P��"�+��u�S�v��㭙,C2՜��|1y�C��l�{zµ�?X�.dǤ��hX��)��B�8UɌH���=B$֋�-זږ��7��b�d�y5���ҵ�� {�줙}�'8��ֽ|�'�_�6��C��\����h��N�z���8~�?��C�/�����L���0W�hxI����Q�3�3}C㍛���&��RM֓ڛoM4�eL��*�p��lx޸sgk�D�lZ�oR˗���C��M{|*�
�v4��@N\��fQ4G��p��߁֛>$�|o=�������(}�$�Q���2�����}np]yյHT�i�ٷ^���qF~�I+�"�Bgy �/�mL�{��!�uO��7&�=���� 8]u?��`�<f>m`�����?��E�R2�wz'��_b27�z߿nq�<��=�;�T�3mQ?��A�LYF�^���:?
(�Mo��L�4�bC���`�Q�i�	8����g0�8�d%�{<�ĘM�#�v�a�<n�{ ^g�������� T׫(<-�dG�+I�Rh"T���-�)B%C�1���֦!�d���D[�������_���,��Y��􀵕0�ыࡱ�Э~�s�_��B����y&�VΔ ���X,��f�����gX�ｪ�[ga��4�م5�HO�-i�E1��j����[���D�����c/���h��t�*ľd�d���z��+�;;�ą��m{3�p	��:8�i��wv�V䓿��K�O��s�H	⍨bP��g'������4��y�"����&V�$�e_�����H��T����և4y�f�n�ۢ� ����3ɘ��j.��o�� ����xK+�
+f����L4O�|�T����y��Ɉ���>�x%���͌A��6���!$E�ѥ�$��ލ=���L�КځۖS���;	1i`��88�KW�ߖawS��j��=^&��NA�i��q~/�����ˋ�{-+�ƛ/X ��D�U�e��!������k���0�5�?�L4ۮ�H�:�'d�՗ds���uݹ��)7'د��C��k���Ց��*�i����\2��zd��P�1MzT�#yޣ�p�i�r�J'�A��Z�]SD��1t�Ł�?t%�������Q n�X�Y��Z߶_�[��\5�ԥ6��<3ɨ�.a�V�+@A����7F[!boL!�ٶB��� ����
:����SuI�v���>�o���Dt?3�7�~���'��t�FŐ��ˉ��fiJ?uɣ0���'�UG-��y�r*y����}��se�����M�ȳ��݄9 ����/_tW ou]� ��fI��,?uI�����Wb���i�`e�l�`(��u=��UO�g�V�4C���k3��N�hl���<#�N�h�i9��=��vH&r�ɒ�17`I�	�,"o#����C���30?��1��G+��+���rm�"�Y�_�Xa�)�yӚ�U��G�Ӊ!?v�c���6*�Q����`�� '���F���0^˩!<�����A�*!��^_��X�� D����r��w#�ݔ�n`4��]�<���(���f�{��[��%ZS�cɝw�ڣ�����|����*_�m�\���o&�i�yc�ٹq��k=��)*�g4�jeɷ�N�6���
�nm��c�z�St�p��w	:��G���q���h�����s�����Ju��F�i'W`��Mխl����:�R�ܬ����ʸI�%����%������8H�S�+T�lߤ���Z3�=7E�1��?����B�ӄ �0�y�ۇ6lj��3���������Nfx��T�%K�>��2Z��1E�_"	(����]����&[�'�R&8є��k���Ó��?Լt�N��p�:&��!�\%n�<�&�`�K����:�F�6P+c�\�oLt;OD���#qNg����RK*�˦�6�@3��3�n���g�}�U�[M���	�PÈWè�'�K�G����<��sUՁ�
�����#���$�i�9Ə;,D���eS�)}_���A�_��Us9��6�+A�Z����-�٥~��G�0�}��ȍ�(��GK�`?|� ������zT��zXXۀ
���|���inL<�V��+6~K+i,�G���i��Χ�r�"
Dc�H���b��G�d@R�?"󉰸1q,�},�1��P�}�&S�҇>ex;q� `G�c��=�[֩�	1�7�Em��e�1y�o+�n'�l�q�4.�fH�c�$�l���FRa�h:I��Ns�:HN��xpj���~�0"�����[��^䱅����Ԯ|lʞ��T�`= ��l�%=:�R�e�l���
���SaÉ����5��k
AP���v�%Ng�7%Hȶ�˓o��|�N�O�� �
�mD�*X��-ӽ�pO���Y__T��9���B/;Z�WU��g&��4�v�Y�ׁǜK��c�-�+�aU��ʍ�n���=�p�����eh�T���7I+,t�n�������ʤ���9YSt�5���x�8o�(�k�����1��o)J��쓊��čܗ<p�Ss��b�
��A9��K&x��-I��\Cw��ZZR>X?�Hjݤ�ծ;�y�a$�#���� ��Ni��Չ�U����x�g)�>�V��Wވ=�AfT[������Y}�?C���3ݧ�%Yo��Ĭ���I��I�1g"�ʑw���3"���>����;yS�����1�*��J�$�1܎�]���U>)����N�Uu�����\.D�#����,b6�6�-8���,2�ho[��������M]6eҋA͔����u+P>y+T3�?k<.��1H�|����%�R����1�*�%#�ʹ�,	�Ǚn"fK��2E60y�\�>k~/���C�e��!�\~�����\}���i+yE9�|9>
(x�����!�߱s-�1�;W��wƸ�z+�8��Ĵ]wZ �G��9C�=6S^�<5S��U�>�@�HO.��V�X��<JD ���|י��}D�ަ�RxϏ������8A|�������'���S�A9��q�2/($%y��VF�]�E��:�d���`Z��4SYɿ9+�>�'ɞ��nƫ�1ll���>q�.�}G�Q��ߥl)����k���̼����n����$��)�xR����P
��VX��G���jE^�ߟ���z����u�T���aYݧ�.��풫1U�����)�(��s��f���������J�������F��m*����õB����XC��kn�����t�ՇG�t��	�)��c���y��0�ZjG�R�oō�����(Sz��=�=�m?'(A󶲈`?���sYjsa.�r�U ���&}��S�otɢ�M��H5u�l���ٯ5�!ř�B�3�r��ɴ[��֘0�Ϳ����P�a��z�=�\�X\V<�;�ẛ�'��Kw	�����r_�X!�"\|�M��	~�ۢ�.��p����5ԃ9���z|��^k)j��u: ���f�R*�;PV� �!�u(���Y�r�_C@O�x����e�5�(X��I�M�E,�N���P�)k"�0�"�ҷŉJ6,�¹��/3��g��s�x������BKqN?��q��!6�q���:��Z��um��!�U%$��F�o� M^�_Ӈ��y��Y�:�c��j��,�p�^*9��V��P
�ʃ�1"�s�- 4B�u�Y�L��ѕƿ_yY�Ve���;A)��
���Q���3�/��#Y��S����G��$�6����&��*49��������Ts%:�K�����r�*�/A*>����.��@)W�.���݇�i���A?���W�Gє�YI�?q6��]�]��hC�ݞ<���f9��$�qH����q��ϊr�4պ����`h�6���{������^��|h����1 ����;��K������<O��c�q��J��k%�Zg���q�!E������/v�b�	AA��p�ȳ�x8v��b�����v0 ���z���V��~��%W����B��,��{~���%l�sC�.1ι�
5��t��" �P�Fxs��`R��&	�gO����Թ<ثΈ$϶i����o�MYl�Ę�i�o��2�zב�c9՗��x�=���Ϟ�Sռ�8��xӾ�Rێ�T�����Vg0n�?�q��~6]��w+��W���\�_u��Ң��?��|��M��~����c�O���㞭ZW�����r�64�N+,�ZaK�r�8������U"���yPG�Y{���U�FE��g��ީUR�w�B'����i0�s8v�/51*T)�`��g����}�����I��y�y�,_٩��3Yaw=W�f�4>6W��~-8�lb1���� (*���CP��k\j��H@��.[�	2�N�(L��_�K��i�C��I�5�����س�jP�6��$���iU3^������"�\�z<F�W�ZT���H+:�'W�p-��H�)Q����Q�����+ BQ��~!k94����� �������=];t%ϞV�]��d��~.K���UmkAq�^K�b$��9�〇|@�����:��
&�q�������k��`%���_�8�֎����QW���2a�2���^��|��~T�j/�P4��/iJ&(:����)Ҵ���o�j>S�q�4^�_��a�x՞�~�'�I��ޏ�T47��L[*8J1%4�@��b i�Q���R� g^4+��9R�5��<%X��ZgT����ΙY�C��
@��_Y�<��x�}�M	,w`�-ʗ���P���gO�bn�{��&F�Y)*g#���c�ٗ����#�{�����>����ב�T�}�������`���"5-k����ǆ	����(�A����&�+B/�<�
(�X�}��Jv6��X\��;�H�������!����������/5�"�n7E_L�� ��;{�_��uo/�E���a�o����(z��������a����M��iKy�S���3���s���c����-e��~���Saʩ�D�g<� �>�u(���%�UO �b���� ږ�@h�w�Y����n���g\.��2<��L6�	�Kx���j_��ރ^���F_���<����c�$c�Mfr����`�g��g���P�ݔ�����D )��B���HV��Fp=m@NS5�d)�M��k�ˬ�%w ;!1|O1x�����Dj�������v�<n ����WI�4�$A%W�$Jof�u�=@�J^�i�^�t�E= �� �������ʇh�.�3$��0K�,Y�
�h���1񘑊�dj�j�D3�n˟ٱ8Qފ�0�ʕ*��p���{��h���3�]4�B�q�wK��M����K������Ƿ�,�~��Z�ǻ Ux�Ro�0'��|¦%R;{�n�=K��I �㗲�aoQ�|@'�#_F���X��[���#aǪõ~>#,%��o�p����-��f�F'}�N_K��X�\E_�7��Bk�t`٘�G�]~9ۙi��.�!F!\@�p�c:I��M�ɩ��;8���H��	��,�r�:�S��Ko��)���'"|@�^Q�A�G���	?��\���X�ȭ�,*�P�)<�}����z5����x�h�=�!���W[N�/n�b_<�= ���)���K�P�&#d�@�WSf�J^t��M{��a3e�>�������S��-O�C�["�`�x��4p�����
Q�
�U��1t�9��g���Z;L}1H��J�oE����l�.��k���]؋7k'��H/�� ��9��5���:��p���;_f����k���W��&,��c��_=k Q�=�$b3:���Xi����o��r��$�v{zs�`G�Vb��E�_�4�7���W���M��ws�^'z��<`�NX�L8��+;ȕ�J5�/gp49ɽ=n�zʺ1jI�,ę�|�� Ð<��.�q���_;+h�H?'QV��WƓeyN��:��G��\k���	%��1Kv2yʔ��Ů/1%H�u��h)�D?��S�f�N]�&!,���{(� 	�>d���nS�^�Σz������Cn:7����\sqꯍ�.�v5�ة�&�Ӡg��d5��}�����b&y��-�=��Y��{���_u`۝���­9��!o�?�P�(5�1	�/��
��Yݏ�Jq�$�WU�N��U�A���X�@�"x�'Be�V͜"������b �2�`��f`Q�6�g�o��sn��*���	xv� �,�Y�[�we��/f���E#�h2q��p�P̟�k�h1W�=[�ڡ�����'���#I�$����s����R�͍�8�XuƷ��3����F���n@-�=��1�?��jp�;&·���q��ư�;{v���5z<�;�K����Z�F��A4�8+��q�)v������^
�zT�h�8�b��y��EKs����i9�6���sQa� �|���>�~���e�ғ���L��ԯ�Ü:X��U,p��|h�(6��n-���,���v^�Yh�@�w��-�}�������|���h����=n��<�X; �����Q�m��1� }Om��{�7���&~�	�)3Z���=�]�o+��W*�?����u� Z������ue�fw���F�u���k�oؑ�4q�mUl��{����Ա�"��ER#Z��M��P'YZ?,��:�bʞVDB��#Js��	�TR�ܦ��-]	(����k��N{U����^�6��0��O#�����X���&8靰ADt���=�cF5$��v�;����-���|;n���xd�����
�2������Ϝ1�����TJ��L�u�����*�e��
�w��f��01���5��I�w���;�u2W�M�F����(&�n���9U�! �[S��h��Xj�=���0fv(�q�v�ԣ�n�m5���Qno�*&��R 0V�A����l��\�/Z��$����B��ⷀ�P���*(.DE��X0�Rr�Ɋ�X��W,hsF��t�麼f#��(C}Es4JЃ�T��ç$Z�t)��(O����Mic��䇮顒�����Q��Z-��	�����P��װ	��9�K����t)��Y�ރ�V��wg��P�ag�h�4���ɻă�Z�R|�?v���Se�C�����$�b�)�9V���?�����i�����g/P'�>��o/-�Y�+�m�ۚ��hD��4�8�>���
�ݥ�h�YB F�	�gәV�T�oq,:N
��b��1�%�ǉ7���e�CK���
������Fla�L�}:����!4_Qĺ��7uQ���ƣ4K CPO�iu�c�$n'@�"��+M���U��'xX4��I-��(�d�ϒ*�����9]"}�XȻ�`3s���
�ã�:Q���B�QY�ǧ�q��|t�xW�4u֢�ŬT��l�R�ޤ7�E=��-��V��.em���"��y�!4���;p+��Ɍ_g����>(Jؑ�پ�_�K簛4_?)�rU ��W�0�[+�o��rJ��`H����f��2�'����+Q�X6z;�F$ �Xf���aa35n��������
�"Y|���肴~V�I��!v��(@=L�l��D�s�Ŋ�ˣD�2VΆwvW�G� �/OJ�agÃb�t;�(?�]� �v�۩�5�؈3B�;@��/�>�� *G)	J%�^^�.��6Q��m� 7:����>m��̛Kq��3 >��󨿩�YV�֣S	^�v�RU�w��9����x7e��b��h�>R���.���C�ӳ�e�3Y��=����V�K�&�6�7/$�\���j���	W8���ͨ*����M����/yQ:KNv�r�W.��&�l����Rzą�=yTN�LV�qܠ��d뛜H5ߴ|'�b�/��Kq�Ʉ�Dya���N�W���ef�{{4Dz��\��[:!�"2��~���N�̖0�/8���Y�hHB���7O�17r�:k�t�� �n@��k�E
�Y�S�/-5:�@8����Ԡ�Vo~�y�C�Jщ���v}i���!�hy{=��"����LW��fx͡�L-���Q�i�GhtV�	��t����ă
�����G���X�Y�O� �Rb�����bk�l��,&b�� �c�`K�˂�qO����a#�ʖ~��W�;/��~�d��牨�O2*���C��$��q���n�_9p<��u���3.�����p@gB_.�h�HI�p�>�Y�W/x��1ky=�-IH���w�E�MA�?f9h�x���0��㥜�gM���O�~��?�'�H����NT��0��ғp���MJ G�â=~N���!�D������b����96OX�=����Ś���G �Z2�9�q���˘=R�}l��!4|[��
[�vX)OZ�}2�J�M-+>���_1�1�ɵ��X$�ڗE�M��p��a"Ȭ��v�զ�z�=&�p;�4��׍r8�\<pƔb��7|O|D�5����5�ҬF�Gq�X���<��2WS��+��x^�ɾs7��@�rv�#�QӘ�X<�x���W�TN��d4�P��I^R���Y.)�/|
��de���Ȯ�f'���ўE�;$��e^�
��w	Ư�8P��)wy��Pi

HU��1��I�`n���Tڼ�⌃���B����e�6'>���7���T*#���+^������Rj��Pb!l��!���d�\a!���g���2��&��Q�b9��v1���Q�[�i�ݳ��x�O&=6[9K�{,6�#��|�d"_�[�}V�,@Vj�Yǥ����^�H�Σ�-r�Z9��ή�p�8v} �^��}�un�ڄ�;��4���D�����z B={�����R�y4�=������/M�@��^�{��th�;�xm���6H��) ��:�}�
��PS����1F�<߲�X74���{R��ṯ 3���r.�Mu�> će��C>Ӗ28����L��zP�à[i_�Z3����9���y��xV�IwA�EB�����o�m��Bt3��U��t";/�/=ưt�N���8�h��v�&�>�A,p�#�mQj�a����i��5M�P�!1|����x3��,3�|�_x�����*E�2F�g��n=��_���fw�\�D�L���7���ӿ�Q��`C7�a�?*\���Yxr0w�H�9 qT��_&q�cūb#�J�i� �j��k�Q@���6BH��3a����h��v���Ѕ���,CL���QMb�ڡ��GaѤ�|����u�G�@�fmmpE~ϥ�ۻo3׀\m�m��©3��w���� �ɟ>*��Qa��������s���<�%OpC^��?�\��r�
��s@��t��%�ݕ��&��4���dʥ�٭	�|�Ѧ��_�'}�&�z?�br�UX>vu�A��k�ԃ�=Zb��K����y�O�n��������t�. �\_�/�5Ɂ�A�s��2f��@�k]�����y	��Pƭ{��"t;��%h�hV`�56����Cr��� 1��G�E֓泮&.e>�0��dX˔:�ԣǂ�`��������zW��L�,��d�k��V~&�U����j�b0kR��=�?�k4t	��d"Rq�;���å��]�i/����K�[��H]�1d?�����YyXm�t�rs��@�FO��t�U�����h+j�Rn{����Mh�I�F��<���<!h#G�-v����8E諤�U}�{5|E��!���)�^?���-b�,I��:��@1�8a�D�wz��&����:-�o��|�H>W3�.�!�6?Ŧ{���w���������ܧ�S��M:�v��@�?O���ûx$9�X���j��A���K���M?�"��o5��ﲿ���p>��bЏ-�g��'��wAȳ�:�Cē�(�&�?���2�GG��?q�i���#}�ҍz��<\��m�1u�+o�ubO^c;�� �Px���C�TZ?[�m�2��"�<0-R��n�3h��ݹ& �ő٢Kb�ܫ���7Ք�M��>�7�>�d,���cj눔�Swٿ㸇"
0>��̎�xۋ+�~5V߳��@4�g}V82&�i'~���xg�Qj��j�aT�A@C��oh���]8��FC)�x7$"],)?V��	�3�i��z�ҾW~WQ��w����/�݉�r����վ����Yө:CwI��Oz���z�W/���)� Ǥ�`M�b���9�+��^��w���-�V�͆FMgÚ�U3�������t��E)��̺(0*d9��8�_{��i7c
ղ9I1�v�@���d��w�	����{�t|�g���!�=���3���tC\���h��!LHQ?tS7�$�~������4�ua]�_�Ȩ�L;��i��9��/C�7'��O"�$f����.F���~^�x�z�~�Th�:1��J��w2�X�ɷ�,?�q~[�����-�\~�R'�[��a�b���}e�2���LKp\�X1�"�.��ַY7�b�v*�Q���zg8�p�"�����B���H���k=�:o~������l���|�1��t��Ʒ��ދq�z�SV<��w,��M\⤗+�\��75t�j4ƻf$�g�N!�վ��A�'�6���p�ó��g�#4�����˧]/��<-��}ag��VFNB������e�Q5M�o��o^f�(@�᛼��w�Dx���y�m�ӱ�Y,�mΞ��M�O��bc�M35�}�S�؟��>�߃��-�˞-�Z�������%��:���ݼF�b2Kp�L�����$�L��z����S2u5�k'��U��yo�"Np�*"�N
+�+ ���J���'�aU�n�f@�1|>�X���������7��t�g��ZVo?��Mh�r�r�;8��<Y �I����v�m[����媴&..e;���N���w�
��!S��c��LC���lzSL��e��q\�}��IԨY��X��N����&2�mk���o�6��
��������i�7���}\�U�Z�]�
�Y�C�>��t����M����%�	[D�6���@�0жdS��iu~g���x�����5��3>)���^7���a���rt&T���Đ���X���2��o���N$�����NS1]�P�f���TH�5����=���R�5��˓��L!H?���f�`��x��Uܘ��0����5�= �=�V���C�*���(� %��/?87�}ypR�j��v���!�:��>�݄;B��E�@�Wn��f!*r/�sۦ�҄\���aκG���g�^��m4eqp|�^?�h�7���8
�O�괜 Uu��,\J�e�o҉4ǩF�s�q�>��l3+û,\֛3�w�	�c���{��n��8�L��O�2�R����z�0ƳSOH�'��%�l����j$�ǲ�r� �Ӷ��ҋ�B����?�AݾB�Ѩsg����7�m;�v�Ĥ��L���c��������fK�yr���}:Y{����@��w�[[�,�Zr�W�>2�B�3�������i�̬,k�{�!V�j��g19 ��ׂ�+��jm�L2�Ӥ��F8a�/9/��dO����i�,bե>�W��a�fw޵��I�fQD�ޜg�19�kSP|$��բE��Yc��4�vJaXw�J��}��"�R��XPP Rօ:=]��
���n}��_W��Ŕl�:��c%h9.W[��z��o�$�:A�s-]�ˌ����2��"'�v?y#��:ᒧS@�1�/��U�ǵq'��iw�M�*���muמ'�ZN��Os�q�l�ڊ��eD�B�[7��Z_U�J�#��R:�ҫ�K���U���3g��dw�!��hq9u�'R�S��{<3l��
���?�M��:��n9�X���撅�Xm�kjL����������҆�$s��{�p�$�����	8�è��F��C���{��8t4�3�ኗS�	�v:�.��!|>W�ՎG�2v�v����OW��dt��|ĉ�2�?�ZM�!������h��h��E")�����T�RZ��Dǉ�yd�#N}�NjA+��<ͷ�3!E��D�t/G����u�\��j��!�B�|09p�N�RԢMn� s;��v������F0���.9X�A�k�>�ӚO�T1U��z0I�cY��J�����ڴW�
�L�s�/7^�#����gK*<�&l��Y;�V����j�5�l#nq���s4��Ǭ8Xl��l.�li	_Mm�eY���n�b���=)�������N���6f�{8nV>����L3$\�?ɢě���YM4���`9�+�x�?%�p���F�tO�#�TU��Ʒ[ˇ���ӟ�&�\[m�� .k$���}[��#��1�l��tfח�Л^��<����.%*�>./��}g-����`҂�Y�-^:���jBiv�顬a󹩡���w��Y�5�\�S�J]j���z�,��1�c�t�SO�L�5ŕ���{/GY�Ry�۳Y�$�)݁�9��Y�fuLbM���Λ���z޺y�pv�L���ѫ>�����%�Y.?��6��ˉ`P��n�I8�6l���>_��˩�p^}�����D)ת�%5��9��!"���Z	,\k՟_c�a��Gsr��m��4��.�L��:򁄪J2��```��v)PtH�S�ʬ;��,?Y<�e�4��LBb�ן���/�s�v�TOtY�	U^����9���eB�ȝ�E{7j�nX�����--����2�{m����e��t\� �A�㹨N�9<K��&��ګ'0�Z�ס�.GY�d`6�*�^ewG��꽷��E�i	��NWܙ}���)��
cA:�
�X-�H/'cd�V;��Q��^�q(WϺ���a]�����@	f<�J�
]�/�MOA�SҦ���>��v?��s�@e(v��������7y�L2*X���k����a��;�n]��b���U$�F���̟~`��|���\jU���?� ��]E���Z�V�M<6����"��h3�iqd��t�"�C��]��*���\x$���	����%���Ͻ��RgL/9@��RK�}Ɵ���]��<�eБN/,�y?.o?v�^����!��Xri����'���,������P.'od���~>2���3��^����Sf���)ǆh.⾝�F:%+��Ye#z�2�sKw��f�8�5�ʷ�C���0X��Y��ʰ	�b��Wb̢	AR����*��y\��!��/eh%�:���v��/%锉hְ$�k+g
C?cεK���7��ϫ�f�ݴ�"�˰00Q�ʐ�sbnQ?�S�D��a1��5� 6B��ӝ��3pi5�u�5f���������f���M��$��@4
(��-%�$���L
��Zj��	�9[��A[��?d�׏^�<�P���E=?A����G!��r�+�,"�865���g�ۢ4�O ��^i@��G�$%Vzyh�OШ���b��l,�RV�1>���,��e@8���s�}�LV��\�S�1�niw���1�����������}#�щkȳ=m��0���9,��8WR�(�s�D+���}���`�+��ȑ��W�����R��z���J�K�Է���H����A�ź��A�Q�*��O:��;�bs�����'��'$�Z�U�%Kų�u�H�ʼ���8�@
�����#�xSjY*y���Kܫ�2	��~.ACR�llޣb��맃w�gO���V�������KC񉪄kD$>��N���N> *�>U����r�%�q�]b���ݣNMM
'#�3��״��u�ژ��R�6��"j '�;��ۃ�ʹ,���m�N͌숶T���o�1*�$C׾���՝�2>ʪt%�|d^z�9C�ya/}4�#WqQ�\�57Oi�U�jP���������W:�J������O��q"�R* �(p:�-�$(��!��ĦIX�'|����g� 9����)�Rjb�s\i):�?� "g?�:�漜��.g�k�����hFw��z6�f1���g���b�nq��zJwXC,�uw*���*��.+�C��3ήǧ�vݲ�x�Hr��q���MrpWY��d���=7�wk�Zxhg?���Z�T�����JH����f�u��_'��8�-���^G8���������a�~+t�>�åP��6C�׾��zp�._9͛����]�7�Hͼ�'��S^P�H�h��#��I�Ƨ�"�M!Y�	�9�s��i;�#&�םҲ~����A~����D�����#��F�o�Av�i���`xP�����^QMuQ(�bJ��T�KU�NB�H�A���4齓��"�k �*-�H	����������g��s��e����gm-����e��{>�w*�U ^��Y,^��}�٧PN�϶<�swg#���d�-��6^�3}���֢��d�j�L"��t��e�uv#:�D��8���x55�#�d�����c_|-��ǘ����q�M���Br��,k,���w��<���m�t�E��^(�_���;*	';�Mll#�m�^E�k��#j��c��DC�Y^C���[J�'�k���O�$�F�u�<�䢣�p��+�4�%ǒ��3�����y���/X�C !|������5������3v��A�	~�gv�q�S�Z#�msט�Y!A�g� ֶ�Y�F$ޭ-�`��T�Z[�۳��8�ޝX#�+wP���"g�BI�-vO���n��m�?b�z9�I�G����bt�ϵ�C�R�"1H̘q���P|{g���1��<�B�Zf
"��#��.f.2�#qh��#�ك�����������o����
�O��ƣ��^�>�����}|x�+��5��%�)JMe��
��{��Euqh��i�ʽ��[B<C}�߄Qi�V���Ҵ���o}��}R)������nŦ��9V����K#��Xe�������\��3��}��,������C37�x�<�1� ��w�Y����$g?A�CeƁ�FB]ܺ�%�~N5�k�#��Շ�/���'��$:ϡW���n\��2�&].�r�<�o� ��ɏs��^���J	/^xL���f���Gk� �3O��߀�E�:�_����{W4�:�"3R�"��5O���C4�����7l���p��2����@��nQӯ\MSc�9�/�d��]%����8��ۢ�j`p�`�E-�ˮ���؀}ld�9�?Ʒ|���;��T[�*r��2�����~$ղ߁�^3s{P�!��n���ZF=V��P�5�q�M{E/��WK���
��I��E��ī?�E`7N�����B����c�^����!u��{���㑰�3�K�#�|��ۓ!�9v��n��<����13r�k�< ��aT?�T�}M��j���T�l�C�^+��E�J�?{�ԃ2�d)/�cmt����:�}���λ���Nz��(�"f+p�v�Ǭ��4h�}�&6R!�1��ۊ}@Uw�s��f���JI�FKcE�6.F�Xۺ�^<��lu��J��;��e�������+u�Z����Pa�
��	�P���>HRTn�(�(sVL[�4����a��Y�l��q� ���:�o��L�t~9�!.K~qD�d�������0� �a��F����{���X�+�/e���(S&�٣r/ڠ]pHd��lw��>#�<Z�_��.�K�h��P�����?�y���`�H��)���/a�H\y8�����l%�,�sW���I�O���[-{z���6�EA� .ܝT�a��wh uN|���v��P�z%��x����1�)@'����<s��\�}}� q��G�20�4��*�Q��X�ME_\�=3�����Sb�>���C6e����4����ќ1�{�/������f��y��F�7�;+��ٹ(���u�|�_�H��vܳО3��Cr6z��=����+u��x>�Ȑ��T�~�'�Өs����DpV4�= ���x��}A���Ρ6��D�qrw����X�t^�o.�h�טm)�X�8���,(�AW�a�q#�Cs�b��Z	E�7���AJRx �g�'�=��<����bE�rKZ'7Lۺ�|�\5��4���6�����%��bPR9�������@�D� ��ȉr����/lrf�8����唖��Ґ�aT��r�%�ұ I��C>>��L��̀ZmN��T���w/�������r�vKS�E!�>m��W@���q�͞������>Sk1�4�A�3�d��ڜ{J����ogD*���X�������S�wj�.h�[��������ۇax��A���f%�I�
�ۛ��	b��ݟ�M�I�Q�w��_r�c��C��/8���3b������~��9�H�)� �^m�̀�K���\"�2�;+LQo�]x�Z?+�@���E n R?w>U\k׉��Z��\�a��ff�Ka��9&&{X]W� �N^����!����4ݘ�%�>�Jb�T͹M(B��]H�3�ɛ|��I϶�BM����O|�$*�g���6�C�� ��gƈ���Y�Q�Pp���]�xD*<%� ��R6�;�s-��UEθ�\Q�B�o�O��8j�<3ݓGXv�g��P߽`,Pt�����NscϬz���<��K�W���C�CI���U��o�v�A-�񛨏}P�X�@v[�̳��^|a-�G�ZKl����M?l�%��$=n.�	��w�D�Nem�`��j�@�7x��>�W�c�Z�X���2.II�IE�Ǟ�U�_r�C��]Vra�&&��'�d��ڕ�E���S�cle��0�M�ҙ:�zq���� �[&>�����;��ej0�(K���k�վ��ۗ�sM�9~�6��ڰ�%fF���fI}y�˴��`��%E����������g��� %�/{<�d��6��S���w,V�'�ɵ�p�Þ�{��@`�f�?��<2y������ct���Ns�ư�t5d'L
l��a$x�Ɣ�*���'\��^�tAb����o�:Ck�X�{2:@,1��_�*pӷ�����"�؇����'�==��0�\ڊW��<
ۭk,�\��	�B���z���6=c\��l��ֈYh�T�[馠��K �j�������V�)ێ"���Ot<����qt�ԙ�,TO/�7ς����Y������oo�!ȟu[u�� \p�4������3b�>F�k�Ac�g��������=�%���<���M����W ��.-tmT��^m?�>���5@=�3���j���z����>����C&��	��:?��=�`����c�����%jp�;6����VI7}E�ϖ�΁H�H��Z�Y��� PU��9�̚r�+���'�3<��N�]v\�G���� �5ۥ�i@v���w�w�� N�� BϬ���<�x�e�Dv�@�>MN�kV>�/�D(h�s��~>���Vi���Z?�x�֢)%���*���|4Gn"SE*�AjzG����ڻ�Y���W5�_u<��>����r�훍�8��u~N����;��8^*�6w(*h�g�t�4@�,%�0k��$����73ոb��Y�Ow09�_�
�@`7��#��%㎯j��h��B�ir��;E�)���$���=�:Vn,�0�?ŷy.�L�?��_L8i��T������%33L�YO::�)�k�^�������k3�N�)���8��^0��^Ӈmc���M�W;�q��摈]+j�g��}��=�{�wKi@��E�L�J��-��6��鯌�X����	A]�������_vpp��k�9�.Om1��|opA�9d&MvPS�u�"̋=S���~��i�<ֹ�vRe���e�}(����0��O虜f�%�&�"ߺ��ĕdm��h������u>�y�K��ۄ��G?I��I��������|�cRf�5r�+�R��L=b	-eEӓ\���^�)?"�ӫgx�Ămr:��v㳔0���b�-o�_�
�������=��w/�C�I��q =�*�L�ʳ�|<2���\?�r2���k���^�	���[�s�Lf��% 'v~�joь�²��H?z�[���7.L�$`
\�����f1���O�W�5�����"��h�麑m�~��3�~��\�f�<���HQ��Й��Lw��V�$�}7$cPD����v�u���&Pn�M�h��Ybh{�ۄh����3$�7�+ж��������mI�����D��_�8h�8��ք�V$�ط��%���0�qY{'��F�U��	2�.��:kƑq"`�]g��i�
�N�ϬڊJ@��5 ۓ�F^WW0�l͔\����Q�Ԇd�����㘺����� �b:/�`%���mns0]��Jz2��ӹ�bgP^Y��9I�\+�]�NG�pL!��Y.��b�t����ڻ�:�]j"䀱O�>h\h<�
P�b���̅�g�������=s[����?:u�2�
���S��X�15D���F�0*���Wf��:ě�>yy]��>581{���%}�>G7���c~�;�������_ �����E�e�̄~�]��yto����x���u�#D�6;ۼ��Pܾ��]�
��~Lλ�Ѳ�1�5tN5�Ǘ"��`�S�*-��\����;i�2���;�R��B�lI�`�z��+���	�s��!{�F�h�9D�(��D5>�Vz�CO�<�${��ā�ւ�a�o�^�$�ߘ����Fs_5�[��`����TP�7,��{���q��$�y��6Z���\���=h#�J� �\�2$uy�&26��Up>�7�+��b@x��}8v��DP�[�tm�����p�3�	b��>�� �t�Y�31�)�a�6�G�{ �<8a5\1��R�D�ѣ�+��}�ힿ��)��p��򮘺T��	ʰ���^rb �ІW�b���>��%o`�`�E������%}�1��A�ԩA�J�Z��	����^�XV�����)@.0r)$��#�aoS9d��� ����l0%�R��B�^�m��(e->>B��A�}[�)#�:@Z�S�1m��Ux[�?s��������{<����I�9~oV9im�l��r�����j�]�Hh^������O��(s6g<^o��[�xҀ^F���Т�fƙ���Af��r�ǃ�~;��
dNu�y�rb�bu���U�T�����Y�}a�>�8���ʓ3Ir��(����Q��8��y�T�� ��t��p�٭����@�j��iS���h��ڒ�l �Y���O0���AJ/���o*���b\�=��S<Ӹ��nd������c�Csq� �'�u���/��f{u9��)�c�}�0�/6�����\�������0Spl�2�4>y'���(0�]��b,�g����I�1��'������u�Eϧ߄��<a����1$¯�2����4�Q7|�_c��.��1Y��/w��ԣng����f�L�\��C�~pcJz}2���_���BL�.%5��5 `Ď�ٖ춱�4r�M>e�����
UZ�� ����'<�����%^
h�����5��`�Zg�:�sP<����zu�p�[Uv ��7�ݫ��� ��p<���S��	��jq"yj��a<G���J� X��۸dd��S�rh�׊W�������#��^��x2�}��B��>�姮J�9����O��R5yH8ly!i47ߴU��(���c�?��]i�S�q����n��?�R^�'��0��{�Ɲ5EH�D��=	/ķ����vCv�� � p��H+�A����kxct��/k��(����|��#��>�[&W����(��`~���gA��BL��|k}�u*J�l�ڋ)ټ'��e�dkD<Bbh�	U�BuZb-��-�ZWG�Y�/�$8�������Ё����1��~y|4��q[�4
��sS�{%p���\*׌ˠ�չ#�a�$���Ȗ\�K����І��ų�A��ꛯ��F|��t����J�-͠��=�Lx#�\�D�w��[����m�a�o}�����W�]��\�mɣf�~y�μ��X}g�"����,�|�`�*�0�[-�a��A���d_��X�;�+V�u�:nbx�� �2�['��d����_F�U�o�EK��#N��>��5Hw��qJdB��:�R3Z*�0�k����푤O��Gڌ��d"c��g��@4��of�>ϊ�28�f�*�:5��S� �F^��Eq���p$Sq�m�4���Y�i�G2,�f�`m��[Ͷ����{�$�v&�GJ�����n�i
c�]���(�|rJ���^e��mL����>���A2�Mr8)�+��iD&G�)J^r�d}�}�C	�t���}F�fB�c��7<��3^�E��k�C;�?�!zSO�"�Avނ�<q�9�Pi����g�@xg��J��R�ӆc�����Z���j?���#̪鸑
9��,��W"�G�2۾��&��b���%��:1&81ئ��q�f&Y��dS��1�Ƭ�!عR�@��|�1������=9��l7��rK I���/K�Y�1԰��r9��a�%R��尥j1��`��8���m,��X���u	M�_����i)�O�x��r�HO~I?������\��da����3=-�=���v��W A�I���N��8�8�����ETjʵ�{��Ɩ��g9m�lx4�8 �ݻZ���w��qߐn�M\�hJt���ޘu�hs��=Z&;?�������`��}�vA5҆}&WTp�Ǭ\θF��������Q+��c���'����x�W�o9]j}��x�����	A1�xx¾fy��yַ�U^��,�܅K�����h׎�z>6&I~(���)�"a��c ʳ�t���10�fn�%.��(��|/�JY��}լ�w9��a$α5A��i��I'����n�8H�<�^�\mc#��Ss�7Z6�E���-�i�P�/m�\h�膟�i���hTʫI/�q�*Q�H;�14�7!8M1_TٸR@DмXϜ��7������æ�e�j���ݙ�/� �Oa��'�:��-g�l�vv����ɀ�ܨ鮱�$2ǃq��	���(�p��\��s;9�4gͽ�:�/6�V��?��+��X�l�@1���e��Yj��iv���:K(,�|ab/7�6Њ������'z�|3��~}�CP���h��k��F��_�����)��>��Ĵ��=`���n�䍾U�
=g��>�%/{r�#����
�a�N�)���n��c]r���HHǥ��0�Ә'���/�#�mߤ��G������`/�F}��1�������}���쩗��ئ�ט��C�i�BΔnP��9o��8-S@�}��4Z3��;�s�K��{T�Rrޑ{�aj񁉥#��Py���I�d�0��d�mo�H-+�%�np�U��,P+��Ԋ��^B�+�/$|��������0��w!8C3�s�79CM/!�nOՒ_���m�����;i�����9_��ˑ��� �6��r�*J�0�ZRa�����TT��?�� o�S��Bz�	=%�n^9�V��Cgڶٜc"��L/C�`���0���"���7~��^�Eu�~e���x�.a�;�~���>�� �mG�]Ǜ;����;%��0���B��X%mw���6�Mfǩ,���L�T��ZiT�G�MbL�Nӯ	)�0�8!����.Zb��?��]�h�!��>��mSXm��1&� [��x��n��, ͥ�&�*y��]�s�P����/sK"����K;�?���af�v9V�Q���=�a�$fnX��d��k}��[��q�c'�9���sV��=̻:[b�\&���ݝZD��&{F���v_�v����-NSɧ=ZzOѣ �_��|66��n�ޟ���l��8
��M w�A����prF����
�a�>�f�Ɩ���Z�;2'��%M��-�x"Y�ݒ����& H�Ew�`��"��Ha>dߏΔ�=p�/T���~��>u��^����[T#"��$@��je�V�7��s�vĊ4����g!��:�4v���`�^����7�| ��6D�Y.���M1��ı�7&��3�ű�kA c�Ƚ>_e�o�eϳ�9+�$�3��3R��,Z����s��/��ǰ9������=�Ƅ��x��]ܼ8���l�ނǅ_�ޏ��xz˶�]
Φ�悯u&�y�@��Cݺ~~�E�x�c�Y��\-�4�_S���b�,�m<����ʳ2�.����h
KL:.�:?%y!7��`}}��T�1�&X��z(�H!vCр��y���=Q� ]j��ܭ&��j:&0�9ss6ޱU��
�;��j�w�(�W�|kBR�<+�^���1{6�&��}�V_ZS�*�pW�/$��]	�ң�Ic���E�C��&Sm�!/(���Fc��Wi&w�̬y i�0N�Bł��.YǓ�jܼ���$B|�G��c�����������B�l�q���v}��� �}�0jM���h����a��~�n�Zs���ŲR����a���z���7%�嚼������ǯm�Sv:������Ę$�Ѩ��ׂ�Ӎ���@�}s1ʷ'gW%ͦ E�o�!4ۏ�(�chyq�c~�����ńS��~��!���kLWa�ʦ�7<h�0�Bk���T&|婒�4�c6��wAE����p���Z�����hOCbM-�w,�����Y��M��'c�T�R�ȵ��V:+��}���NƳ�I'b�0��o�ĳC|�E~�1��g�dJ�P�-��{�UHj���g�b��l�1~�Q�Z�N�ѣJ�f���ĳK�??t�&�	F�����������>�f���-�E�J�xk_5�����*���ۙ�y���Gc��dꓼ��~�+/)X�E���E��zІ�k����!��ZgWML��@�{?;Q����P'�'8R�y%��S�t��Nϗ�2+�c6ڒ��-Wa ��V���W���VR	�@��_FB^�I�)�W���A���T��!��\�rquE�GiCT���r@�O��V�ƺl������Br*��1[�*q�=	���tN�c��)y˩W�,',�}�����J&�����������o��
�M)��P%��䈣#*f�}Fn꧎5��15j�����lwFHb��'m�a�RA��cI�\�Ã��Q�/ܮ���c�u�9ב�ݾ"��͕[�����&�S<B���m�k�zy:�B�GE/1�u.�4��K��I�
B���K6�q���.t�ƛ{Tjf��e���Xج�<qz��pײq@�[p��~	 49T�XԑLa�x;O��h�r�D�9���hO+�7Iv��րjL ~�ë4��ƥϋ[��ǵ�
W��y92gm�b
��W �髢A�u�Q��8c��5�
��@)����/e�F��ۛAw�A;o�`9����]
0�џ��5G��v(-�������ʆ�%��+-eŊ���6<�#_2���D7W��*��_(�~�nGX���&;+3�I���S������*/�^M��/KAn_�����"��v�9��>i�G��0�
eg>VpL�����O�v|�"̒-w )�����\�਺�J}�t�Y���՛������N=A����2�8�z0?oꤎL`8�kjR���R����A��6B��Nӷ$o?�m����N3��=�ӂdu_o��$�W#V���f������J##�4����V�9}��9^ZA�{���ɟ���%S�T�˭��Ll��vN��b p��L����d�-��0� ��Co��������ZK�ѳ9�����4�Ҍ[�};��[��?~=�aO��k��8e�k�y �A�[fY@�VCxH��^��O�%�� ����̲�"�z*�XK���wи�1049Y�`@�|��ބ<	僌��E�" ��'g���&�n�*���v�G �ϗ��C)�W��ĔL��g�냫m���%T$��8`�{�ῧ?�5������Vֿ����<��r�A�̖�T
�Ә���W����s�%x�������B86�Ti�H��9���u�|�X�/ɸ�/85<���ri�8�%a����ٗ7�m����p�I6A_���r��>s��	3�'�>�m������� ��I���W���!���~c��^��nE-fȜ�����}��NEJ�xf�^��ޒ%<\����џ����L-�S7_z�3�Ȥ*�;^~�������>�ż6�k�F�Z��\��(F&
�������'�5�Dj ܲulN��	Iky&9J|�k���S
OH"����A�IZټD[g�x���C����_��Qq`�p^�\�����j�6	"~B��C����SvުԕA�H��X�AbF�<�����A2�����u>w�Kݛ�Q���}C�e�����,�}𡉙�ǴNS����R�
��`�lj�W��s�yx���s����qJ��zx�]AC�D����fԭ ��4�(ȉ~+����zn&�
$C��0�� _xT��A�ז3�9�n��Fk��U�&����<�z$x�T8����T��8�oZ��}��-��Ȯ{�E%K{j��G0>��+������Dԩ�BYO(�ئTϣs1�38Ȳ=���\x���5��ў�W�	�o7�P�#1��X�0Y�C��uG��|� o�<�_%����ܕ���A��뮟��o��7�[�9����>���6��҈����'3�>��/u@�U,:����$�"?�Ժ`-��s�Ee�$��g�8�i��?�m3u����a@�����|i��`�*�����7��� �]����x8���;	E��Y��*�M�Y

<�d7	��@ni04��ǀ�|�����r�{|��rwU����v��wӴ�s�ev�̖������L��8�"�2�l-�����E#?��D��e�ԍ��=�6��N��W
}�Tq����Ώl�g��=Z1L���x�����R=�"@eeͪ�d����u^ud�2�Pp>D�,�A�0\%��E����(;�F-�����l�L�hg�6x��T��m7ә{��4������Ɋl�}����)��7��2��&ӳۧ���|�=�B4����%�h������ӫ+��zf	ˋq�}n�P;��=}m��8�s���	�
S�2MA������`3�$�Zq���;�y����F�ۊ�"V��ۍ?~,QZa>�vZHn���{�$kǼ�GV���@vW"�h'�����K�#�g��i9h��!��`A�bE�Zج��M	{�o;L�����-�sإ���*oq��/'i�}��*�����up����I*K[.C��Y��=r~��+�R F��q5�/�� �S���	>{��Ζ �K��ܽˎ�5,5.o��"})�v,�@�c��D�;.qA�A�vɟۥ灟iTv���q��,���V�l>��/������_|/^�
����#tI��	�lV�B�g���s�6/�F�]_�w�Is@vx\��6�g�*���++o�vl9>���\�F�9�HM�;��Ѓ %��O�<=�{.\B� �.`d0����|�H����H�8���6��[(Ռpv8�$U����,���҄�G���%�뽑�s�����\�<1{}D{P�R~>�zb�[&��߶�@��l73(��� ��Rw�'����~����"X���_W	V3�zaF8@}8�kkrxP�k�t^ً8ي�fA?Ǎ������Q�;����0��D�>6�b�ad�>M�k����L��)Sʻ���1��P��_�+�؛��쑸���D���{^Vd��Yʼm�½�v��*�R�q[�,�%��.��92��i��脺��ک�q)<�<T j�}��ۤM�O���������r�q7����Jg���8H�g���"���YZ��z�<ߍ��}�T���0���%+e�T��nc�/`��#��MɃ7GO�$k�=f\��Mh�ӧi2/��:��7�)i�9;�g�1��ںQ�'�A�̓�j�m�Q�3AzF����Z��l�B��g���٣�E�Բ�7�F�U�~���Yo��H���{g_�/G۳oYT���uz3�J$y���l��X�GQ�y�4�)±9s��`���N�����ۣ���~+�\��U���0�����%���ԧ��A�i���!!��L�Yi�)~���gB�L��������JފbEM�7�Eǯ�Y��|�\c���1�ӝ��\g�
K��>��y
� U��$Xae�Ol(`���"��퀈q�z���m�T"5/4�<���_ҚLٸ-�m��;�J ���&VL|�!}3h�������V��U3[3��,WЯ����sk�1h��J ��D&��=�E[!��^:�u.�ɛ�\@�|C�%Я�Պ�+��qbv��J�v�Φ���zɂE�Yʊ�Y�o�t�f�|�h|T^Vg��w.f�p��K[���p�kw��u*
e&lr�F��KDa�p�|hn�\�1M}љ�����P�;�����Յ������M�����Y[���̂�i��7ˡ問�h}g��}�f�`�&����1�T�91�84�=�|<mgd��ٕ�����}E�yw���kI�	�XB��+�u����	g��؋ 6N�~D�6&��p�BC��\�����5s���$�
���O��H��R��䌪�K�i��~��4C�.*�a�5�"�@����#�����@��h�8��Rw54!$e��w�%<��s�4=��"@p��Ǥ�D�Ahra�p:G��]$�a~3)��K���N��
�δ���4��d�i��Y�ք�݂^(����nK�]���ӇXRM�}h������Tf%�E=<*a�����N�X�~�7����7�uY��s�{lo%��ߍ�����y�;ڣ1}}D��Z���e��t��1`^h���KE(�_�On��������FQI����
=������	�Iın�\�����/�|p������9mQ	�ն�
I	��u��T���O��D�k�zW�S���6�$.���C6J�������}�A�t��㦣�3�R�yN���Rv�\��'������Z�gJ��`�
�ْ�G0�����NP�nO}����-j�w�a�<5bȸ	:AGg�����m4mƽ:(��E���t�. R }�lL��`�濅~I� 76�$��:�W4����X{��;r��8���&k���v�y=_�[ٮ��`n>���'��5t�>�3��h�"#�y1���-(-�k;���B!�/U=0�26���X����o����3��G�)k�s��zl�P�x׭�z�=�7�����&��/
��(�b����dĪ�ʄ�Gu�.�����
�q�^*뚚n�+�����w�	�4���K鵽��#|�F�x�՚���A�K�ѡ�&g���j#�:����VW���U����r�F�b��k�N��Y���t�D�r"$��J�OTȪr f��%?�bB)o�"/��`��$сp���+�6�˷9��L���D�)S�iݷ��Hk@�
�E�TO��y���'�}
��n�R�$�KW.~�y�
�:���3R��:&�� �;/:�@}���8.��P^R�|��1VqN]�>����g�=�v�d�����1��TL�=rYm<]���XS�F`��l�V7���^i��I���	�Nܻۡ���wen�xn����,�/�693�<�h����&r�s&��Y2���-��ivl�ƞ5���[����C���������X݂�${M���F#,��e�u���vz��e��/+�N���&�ŀ4�Y@��P|tr�v�V��\�����P��q�	2*�^	Wm�i2�^ë�:OQ5�E��ݳ�:V�V�kI��G"��)�`?����� �6�����ꭋs�H:�[ޅ�F8�\ A!��}]����I�c�Q�#.��t��h�Z�������@���{q<�=�?�]���/�^v�i+|t�3u��*>F�V����N��?��3)ţk������������k��K�[
K��(���-�@|e����g�q��I�s�К�㡍lV���'�t�K�d��2��JJ���?�5�GU-g�^�D�n$ɭ�m���;����+���{��w
�k ��n�����$����h��]6		��'1�n�t��#��1[>h����pdA�=�Y9�H��\�M��f��$�G"�g$a��>�(�!'�f�P�f�|O'L���<fC����e��,
�k9<	��чڛƸ�A��{.����8dW�)?Q(���~>}$f�����ϐcmr����VxJ~� 	ݰ�H��_�қ�|R%yq鿡�_�t�2pi�z�C+�}kP(�U��A����z��r'�9��-a(4>����0^��eϷe�����QbL�H�5EϠ���ǖ|�6����=~~�	|/�fC��kE)0ߵ}9v��h7٦�]��۝fZ� s}��n�}�reZJ����ZЫ�-n)+E=���#f ��	(���_�Ta;����5���3rҕ#}+�/`�A�se��,݋���\�愃�э�����h��&�7"Rh|�}����Cx�z7GK>�#	�<�B�5�������VnIG��o\��^]^�N�Hp�Gu1�˂D��|~}]�cI��g�$��b�E�*ɯ��:%���Q�C�NP��D�g�0WϣK�����!%��koK� 5��Xa~�N���E�m���x����Xӿ����$o��A���wT}M��jAt��Dm�G���p����0Ug���T������`l��ۦ��q5|.&�3�,��S?e�Ҝ1Y3�������xL\�
˹���7u5^1,J%�ڎ�,ڭR��n��|MpQ3U�}M��e�K߈�%��A�:e5���\��V�s^�W�I��X�<d�O��#eo�,⫓q~s�� �˞3Q%����/L� ��'t� '�I�@�x��_y$���%�rg&�U�|ɸ�<�I�w+frD��3Q��D���&g���ǜY6�j�ߟN����.��w�6?�\���e�4��7�˹�<r��h����2���ʗ�����~�Cbp�&�rp��S�Ӫ�t�<��|�(T*ԝ���CR�rRޭfw�M
?4ѝH��M$&��0��9�ҨuPp�אK3o؍�D������J�k�]�pkz�u��Jq:�L[��\f^O�OE��&a���j��%����C�g��B���XUa��:�}3b�|k�Ŏ6ݡ�5�k���)Q��|�["v@��� (�2��	��K������wl�Mc�B�+�?6[�鏿�~J��g`H�.}��ǧ��b4�	ɹ�z�Dw`=�����֬a�,(�8P�8;��Y�:Ÿ<�,�4%.�r�Zc@��{;js�B�����3-e�F�ˎ���[�
/ (�螰N�Q�vv�����|�MI:��QE�V���Q)M��/�2ZI����r����Е5����m�8��I::�q��bb&�o= 0X��?�n��x@�r��qSL�<vi����ݐM���?rǪe>��{���hCG']tyZn�TQe���y|���urD��G#�Nt�j����~��A������I�}U��m*���,t4��T�������5K$�`1��^�������d?�K6�ǿ����#6�Ӱ-�CN�4���p��%$�CT�B���_L���{�14�H@�>�x����_�܎�Gk�;�P��Mp�8O������r|P���nc��S2�)m���?ױ���jS^7Iz�M�Y4{lI��v��ڈϫF)w"�qe[��߇t�_��&UH����k{�aC����D ZйLz��˩L\��@9����_����F�'��x��«�\�q���tt����o�2;��xawvge��h��R��m�5n��/q<RI�i�ߵ9��KKx��S��~�����?q���~X��e~8;����-7�y��1��?����~c�raه{1`ɓ��N����i��AG/'؍���3���]|��.�S��*���!���hT����켛z��_K�i_��o�2�ss�t���T> f������Q�ng���m_����n�s�3�=t������������~ +��l_�f��wV��(�#���N�<�&S���;:�Lw����y���P�
$��`.X��S����[�W�ׅ�˜��_J@-&�p|���~����=T��Ѫ����wD�ʭ��oD��<��_&��X,]���;=�������.>�~F�|���n����k'��<.���u��7	&V�:����Q\���5�6'v�U>�G� �SG'��m��+3)�	�搓����<|D�~TtF���GB�nk0}�,[�a�)��l�������t7.�_����L֘ �ԇ���a�"E���d�3s(�7 �`���K[�sjsy�d�h�w�|������5~t���4;Hz��X���y��1��H^����ƚvB���L��ݵ�3��{�.#|�z�so~W����"/�<u�7��wyd3L�ƞ6�#��M� ��� ��U��b8=���s�o��{'�����/ ��C'G�t������&~����cv�3��Կ�Q4�(��q��� ����}Sv�;-�t=� @�w�k��A�Ѩ����!/l�$#��;��O}��;Uб,��մ5F���5�%��,���N֗�	(�?�~�F=!�>j��{��h�[+����'ϕG{���ty�s�M0{��=��0J�ȬYGo����Y@h����5!�&�.�=�h+��x����r뵥	�$I�M�ʤP:��5�#y'o0��~~~�"Ndj��ȯ���*�(���|B�qNa����'�	�:*8�p���րA���g���R�D�d��ۻn��Z�9$�-���M,���HB�2OFB2_H�Y]�����\�zݍ6��uJ���A��K2��>�Rr^]�6."�@�TB�u���/4~�$·�a�!�;~T�@7��0X�m̷>�n> ��7p,U���A���,�9���umw�eMAA`��oi*���x�]��:�D'�pk^����pJ@��������'exj�ܰ��Z`D�WܒOe�9�������-�_.k���/xYH�ǫ5�W���W�y����1b���/�����I����C�[�5����C�Mp�(""%���%%�1b�(�Ғ����1)�́�h��=?�߃��������]q��+�����t���O�ڵ
�I������"N�u ���g)~لT�p����t�?�������H���~�{n�V�%�v�/�Ѣ�o�R��=����`5�s-�Z�X�=C|o�2�������0�X�<Y|�(Z���#�z��_K�듳Y�0��k��vc�1�&v�5����bTo�V7�M}�Q���<WH$��0�)MO���2ˎa�C��i�@ @�����]oJ�G@6�7�S���Q��)HvZN�GҦ/����Z��q�⣭O'>��,���{fJV��e���iXQ��Q���f^�h�*P�&�ʔf�%���Ew�y Eew��h�	�ؔ{��i��VK:"a7�.`�B=fpcN���i-�*'S�����Ӣ1���\����Yed\�P�'��<�"���k|��葼伐A�B�\*��Y������鬕^[�+�����K���h�5�$��9��(x%����`OQ��*A�L.�I(7U�RC���ͨ��m�|�~Pdߤ{b���`� ��"�t��r�~��8� z$eK��R݅]@�x�K�@���)��	������ɰ��VxGCP3m�ʹ����̍�j�Vl��|�c�W=&U&-����Mb�eG.`�EY����T$4����R���۱���7���_�-r~}t���:�hUa�j�K�{��3үX!UE�0�^���u���]��r� >E��~��P��0C���a��f����5��]�����i���K�����C�����(g��ܕ�y�{i=�@�;��[}��á��!g�1�u�(Io	�>?f�e�����?$:/�,3(er�(R���p[��+ �%vv8��	t��s ��~5����c'�o���@r�x�%ŁL�ϼ��p�&�f�^��]�M���e��d��ɕ1����<yҟšZ2FzC@`��TZP�]'�9"P@d�������"k� B����I���M�=��pn B�A���~�<f�m�G��{u;0���LܰD}������+��ɖ�-�Z?}�4e��:Ô3����J��1?�a���իtqw���p�+�k�8�R�z�o�KIʆ@9R�"6_v/ ��0�|[Ŭ�ʾ .��]���s�/A��7�H�o{~ΐy�2�|�.�i �l�
e5)Z��Θ��6�j�!U��,�*t({�D3N�/v�C�]�Xv?�V`� ������q�������`�jlQ<�SB���ayV3�c���bP N��DS	���Ad��4�܏8����5"��S��"��s@n٣�)�/��	u����%3�o��Ğ\�ޙ��-�t �?i!`J�,��t
��ʨ�Mb=bF��Ŝ���u�|J!�_!v�C�K�~���[�kDw��usW�����"��ċ���mG�w� ��۴��F˩��-|���B_��A.�� =�8TP��Ҋ�w��3�Xz�Jo��!��:�_�u2W��p����O�4���B
x����G��c|��Q������sD�e�U䭑R$�'��%>]�|����j;Bs�X�궫��"�X0��v�Ӈ_����{~�3�-?��CxQ�FE��>��o|���q�ݬ{R� �Ă�$�TI�ˢ]߀���t1X�z�$�M�jVl;fN`�<��Q�<����08�8n@E5�����DBm����o�ɢP�s�#5���e1��m�%٭:y�Kդ
P�ݩ�W?[a P8P��%�>1�c�` �)��Ԁ�}�:��ta��{#��7 ڡ�oR�ղ�|�H�R�g\�B�_X� ԣ�5`R7���4+�?��o�ʸ��:W7F�v|li�	��q}Ơ��)�]+�*XO*2j+m�G�@>��F�H=���v�i�Г�$�Skn<�)^�u���i��S�8�'#�2�A��Vꥅ����L�V@��b�m�6)3j��d�_w���e=�����*\'e£��,)h=�1ۋ��Q��9+(�y�*�~�TS�ͪ��ߺ&��n	H�`�k�B��1�[�q4�r����C�s��2��σO�%'ruzB�����c��4 v����R��ZC��Y���l���);̢!�a�	c�����Uy�(+|�L����x)b}�h,2���C���\IL���[(�����z���3�q@R�;��S�2g8����tW���H�t���"���~E����Pf���s
@π7\ �"�&7�Pk��N�o&��F���x��@��}��8^Gh+��g~�%'�����O�a<��fB��*��~1ً]��m��JY=EW>��F�����ߜ����l+�:���0k�y�P���9�FL|ڸ1��.�.�N�Y�4
׉�8�:�};j1�J�ܘ��?�[;�ҭ��U�7+��/G�<�W��6�x(��ǥ����4�!�ϋ­���L�}f�-����	���<V�y+�'i����B��ih2���E��7S�g��
%4�S���04�Զ/����]�Fԡ�i��Β�ɧ��ԢK7o^�޺�7A�s�ņ�j�Y<�<�Ů3�� ��m݅�_ώ���K��Ee�"��o�m���zX���]�&�;��S͵�[�ch�Ä�s9��f����P�xY�{�I�u�g?�l4�&����)X%����6-��i� p�mWF�z�{��XU)���ouM@�p��8)��,	�4v��,���u7̵�&�&��� ���)��Ar(��(U6\�5_I��,� ��b�iԉ��psx�S�Q4X�Ӌ�A�)�xx�H���S���ҪAomI_��s���l/�oo�N�)����\Jj᦯v����E�ޞ�)N�Av(���~#y��O�ʶ;vb�u�^�W�f���ĞCG�!~�#��B<4o՚LZ���$j��loDVb���V�l;����`�3\\�i���ea���d��d�rF�^2@��xx���<^�=�h��,>�*^�&B� �60x7>`��Ӷ�A&qx�p�i�#���jt�V#N�b���H��/^u�h�ʁ���F����w�<2McO)�E��&ZoNI℠��
i`AA-�%	�p.=�'��b�a7�h�
���S?�&����:;��� 	$lw���`"�F���O)?�<��cއ^`t4�.��	>�D����oY|�M��3r��g�nɭ�g��\�/�N� tw�袱Ǯ���*cFYD�PF;��s�D�����%��U`�b"���=z��4��P��w���)I�lU�{��J[���ZN�>��\��5�F5#;(R�O��las%�N�c.@d$5'F����D�Uu���ԛgǧ	��}R�-(�6:����H�`�6D�rYU�:�htk��,�{�P�3d�`�-�ۈ"�J�%���օB=8y)�)�<T�����,(b'����{���ҍ+5���	���l�g��	��K�T���� �l0�n��V����}�ζ͘OY�G���n��:�ZT3�U��I�_�Ѓy��G�_�fC�*�J�sT�0/*#|�V�����6z\����|>s�`5��.�.����f�O�ՠ��*R��P�!�l�m��/O����
`��I�D���.F\8����uA�v"������Y�$*Rx�"�Rq9� p�g��k�"Mo���1E�~5c�l�s��-2��i26�Y���r �u���-α b�l���{�G��d�E��ʝ�γ�#[U�x�S`�D�� [�)<�vT�}{�j�������wRc�8X�l�_p6�u�/:W��|�CM��U�G��	ՆL�����iع�c�V�e�R�tS�����1��m"�ɫfT�w7]ߚM�❡�h��@<�w	Ke'��5�vC�&N`R�@l�f$.�]KFe��%�jX��;�&0���L�\G ��L�vE��Z��.�{Hk��q���v8�فh4��&%]�w,З8w�ݪj�[�sj�a�Ytl�5&YY��8o?7���d^�.f��g�&3�$H�RQQc����������ܢB�#�P���bL�� |�5]�V��Ϩ��
�C�x����9j^4��cLM��ȋV�9I��g�q]�K)��Iu�w�4^w6���F+j��f�����*X{L>E�DY��N%5���Z�V���B�8��=�vJ�[���-���S�T~�N�[��3;�+[���`S(sC�j�'1���QLKzw�f��"�����a%�W^��#M�Ǿ�S��mH��,]��~���>�;a�1�q�o�	��D�F8)�%+H)�|g��* �A~�l �6��а�g��tn.U{釴, .�0�j
��@�U�K�ɂ�D�w+�.��	ݺ�����o��{^!4�O��Gފʰ�@RݭĻ8C(��N�����L�ʚU
�J�)\�q�9)d*z������p��
X�<�2z[�s@z�U�Ob���Gf�Q��O�ᳬ����j@:�wn��﯈.�͒ݏ/�ͷ�*�ڠZ��y�T��ޤ0�/���%�!d�Ν�7�tZ؀{@�Bi[bUP���o�������  ;��l\���W�
�ïj�ɍ�f�剟9��G��PB��>�:@5Ǒޚ+���@���0�).o��-Pm��ֱc|���.�1��312~��o�z  窂S�d�oT�I�J]�Fn}Eu��U5���qvwj?��9Q`&��1���������%��ɭ+��P��<�'�<��
$�0�{��_�KW�ք3�|s��F�T�W�ݐl�d�n/
���~<K��!���V�N!�YH'���Z3�e/��PiY��U�� ^�����!�r8��w#�c�(x���|=D�h���iJ��^��м*m�qC�Z�e��[���o�N��k��d���^]�d�c�����8�ӌq�P�C���r���}��gV#ecAד��V�?�{S�e�+�yo�Y���y<�j_�%��y��#�Pޘ�[}�
�Ƌ���-*�+����)�s�׿�H���Î����UAc�3�T`���X4/���zH��+?AW���� �0�
jDI�&�
����\
�!����߹�B1�{��0t8`n~�i<g�(��U�n%����3�� `>^�4��]>'� :s1PU$�ҫc�qb����F�)�vm1�{ ���U�t6;�h��D�8(� X6�Y���#{;�l�a�L<� t�2S~�M#�@R$�*�S��[��+%ܷ����r�{QI�FS�� h�H��j��/T�yQk������]����!�~��-O�(��a�)�,����&�B�b@:J�u�#>�-�K�������uۥ:��l��M5�:�W����f0%Әf�����=w�$�� #�#���V/��263�~ �����6Q�N��Y����� e���Es�b�Z�0���EXVUѣ���wv>s 8<�Z�N6	E�n��7�]�Tj6rO\�.�lP��s7��׼����K�Wb'�sa�sX��@�W7Uw P�Ve�W\�w�=G��(�x ��c\�d��:���Km����;[16��y�4��8}����G�Sk:�zk�v�6�����C�ĩ��9�@��\p"�1Dс�`�;�|����-&[۞�[...{�
@�L������gU������ ��<�Tle�Q�|:~�>�t��?g1>?B�j�L\��e��sK�1���\�S�G��������I1w���G��.���I�YkP�5�P0l�?B��9��Hki�h Ӹ�TT�o�hXJ�zH&���#���a7ŉp�n�s0�x��0��e�����-y�b@��e�
�sV���]to�}�}8\��+r"Ǐ��>�ip�&�꛺��V�
�F0�&�����E��A+�_
�`d��(��[����Q%�u؞k�A�&"�e�4]:���pW�i�x���y��Q s9c�U�@pU0$�����%=�9P�X���
�"C
�D!�����qd�>k�$�i�Ѱϻ[�b4=�˸��<�:s%�fe �vo/-��cI���kfrS���1�N?�$ͫ��[�[�Z��QJ@Q�E���w3֍8(��~�FlV
�ɮ��b�򶑜X�q�U�%��K������ɰ�(-,A�� 5h��(NʢoQ��p��{��p���+��Rp]h:��.����Hl�b��N�~������ӹǬ={`�Q��ZJ�?E�X�6�hB�)7�3�cb���= F欇
��~�9=���KhU�k�(6��Ch1�w��M� �ǀd뛏 �:�
�|�2|q~�^Q����"���6�ulK��Xа��DZ��RBjP��Gو)U��'������p�(AL�"R�S}������m)`{ NP�0���|{��B����Q>�=��ߴ9r�o5�~gx.H�)�S�T,Y�����?0l�X�{�} ���wh�ʄ���n��ą9 G��=xC8��Sv�p[����v��1c�w�_��.�^�4���M���P��z��T�'e�'��g(���x�x��@��~���V'��q��3��K���,rAu@Ej�2���]����{s��3>���anѴ��"�p��k%�A�R�&���p�?��~��� �T�q�Ƿ}v�c��m*Zb�E|��d��*���8.���׻�Ыr���i[U;���347Qv�|V�Y��B[������dG���\q��pVfNy��R8����C�ț;�ߙ�-ٵw$�.�x��F�I��M.��Q^����v�J��n����Q��\��n�;#s�6Nɳ��b���ٍ��(��i'�{p˙)�t/����Aq�e�6�!�M�b8�0 �.nSݛ�H�N�ewl�Ǟ��s;���(��� ����g�U�&�6���H����6�`�k`A;Ŗ�.�=��na��*c�T��9��V%�������Ұ�g����"�d���b4h�y�ة�M�9z�Y �9��|A�| I���G@�����:,wˠ~cCg��ޯI��=��o�NU��Ud�������>Cy�kFݸT���4�?��F[��qÅ+��� 8�gv*ix4�n��s��(�wX)G�^\��-��Mu�S�0��4ai��A��r�86�^t��v����;$�	�Ir&�����6=sH�+���4 ;�c�:z�)XRhg����`}��PR���1e��gފ'���;���h> ۘ�}��af��Ј��6�U.UC���*I�yJ
"���<���2_�G�q]FH�28BP��^�T���i��Q����ʒb�]G�-A���\�;���]0�� �A 6�����!�ۅv�JZjrt���*�kJT�4��Zu�Gʴy#۸�%����"-�����NW��*~heh�i*�?~��q��6�N)u��Q�$�u����׿u�*%��j�J��a7��X#�����i�M8)��T�.K����n�u1�gƟ��VAQF���� ��8Zp�{�h�'Z/��C��������{����q�����P@f�Y�1SVÚa��L:��ss��<��VP.z�X�^�x�?k�p�&m9�4#�'�M�P�"	��D�SMK�[��J�2���g�-�(��3:���y^��O���\G������w������������y��c��Q�����o*+|��.�t�3�e��i��6&�q�'��Q�N��c��:�`̵�X��#�����.ٟ�g��1~\#��@��@�$,ä�w����=��^��.�<��ɕ#)��W���с�S�/����}s�/,s)�D[c�dM�<��W����P��ӯ�������Kk������V��٦���y�{i�x�[��m$�A�b�@�G��<&^�e�1�ˆ����J@�%	X�/»�\���!��d{��=�v^m��c�j��/L'�j��Ώy�k[z�~��Y�_/�4B+n��e�u��Ҽ�W�ƷL3�9%��/V�2k�#)^���}lr��4�c~�z�fH�֌��ˊ�I��\�#��B�ܿ.�����������.�gB�留��@l ��L���P���=�R"�;���ww��4җ��
�~�#�]���~�̭߉g��ݪ���0��)AA�� ��'���^��BAb6��D:�����n&�l�^6G�6}�v�_~��E��@M�psX۵�W�a���8��ߝ��c��q"M��H{x
l�]|�v��f0��k�(w��IzV�踏:�<�\#%����:����x+h��jC�"C���hd:   r�yU��4�.D��K�W�n�U������W��g?�k �
�w �GĨL��&�Z
��_\d��qg�͙5�ʡ&mr�����ҏ�)1��œq��푇� V(�c����5%�1����972r�+���(���=�kQ&h�"=���ߝ׋���XK����%�o ����s�bM�ܤ����,R�f�����������L����T��+�f����u�?9�(/�-����?�f��?^Ky�M�;"q=A߈����t��2p(���'���7�qu����~*��x��I6r�(�fF�4�-��9A��y6���~o�9R��Q��<��n��n+<��6�%�t�}�F���A�I��
h������7����������P��i���TR%^�E񛰺whWW	��T;���_9!Z+gr�vs#FEV���m�jF4�� Q�&D�D�F�Z*�I��^d���#�i�	�C�\���Y��͜���&��qIȃ��#ٕ(>���қ=p{C�~1����[�қ����Z�+}[����M�ʇ�磺��xbr�Q�$�PWۉ���]{/$��_�<u�X�a��%��|���2����������Zv�Gy����ZW����.ap<��o�:�U�4�Ϗ�P�UT�a�:��T{fh�#A�w}
%
���P?m��my��7�Ct�X7zv�!�nb����m�@r�=��a�����݃����_+29�5��+��*����;m3v��k�\қ��=?>��/=j��T���5B$|	K�8ف��X<��M�hJo�H�7m��=Z����T�������h����ު��h���9lw�=.��@�3��?�����D�z�:Z�}�tݧ���@5��eN������^䋴�3��ہr`��yF�5%��ٲ>��7%&��$x��M�6'�lHz�h�{�n�ɽHUe�y�>���4�����"��g�*�����׈��!%.~� �}~��d$xL�>��,u�n���)y��f*�#��Zp������~d��J�>&��7�lMt&
;M����7�Tۼ[�����ť��4�@��Y>�`Q�/��/��#�-�n�}׳.Y��)z�E���qj��N�9��.��ؖQ���}7�m*;��Y h��;Q/��m{K�l�g�����޳R���c�	�d�F���d��I-%�����W�6|���-���M�90���S|k����S���g)��;�c�o�!Cb�П����!���E�$���=�f_�?���		�<w'$���7Iț��]ܮ�i6a�i<�Z=wky�6��x��BW<�%<z�����}�pe��� Pn��C�z,z��)o�<������+�����dc:�aj�K�AW���C����N���Q�g�mc`���,����G5�
:MO^G%'�)��F?Pt�?�'�����@|M��[�W�ժ��$Y����#�R-���Y�m��02}����S8�m��5��s�r�J��K"I� {���Ǆ�S�[�Z5�����a��%�[+��3a��lɿrT���c	�F�d�ΤU�#M�<�����n�����_-�� �b��HDTP���W���mJ�tkV��Z66:�B��\խ#
,E�Q�p4�y�i��x��L�Q&Q����Do�!z���~�E���+�D�Wv3�yϧ�N1�)�W)�x���Щ�)��T��,�*R��"e���γE�=�>-Ւ{��p�; �=x14Q�n���lqY�N]kF1
^�w {�R�M�'<&�}O�t��bF�M�l�W0D�(�]�`�j�����H�� �N�%:��
�19H6]՟�@c�b������H?�h��EW�|�"w[O+��=@ Q22�F�����k'�q��:_�(Ķ����7M1�y�n�_��:{���L��d��/�R��O��ف�Z���{��^XU-B�a;�'l
���9���A�4R>`@{+깞��q.�'�w��{e�\ؼp�t�+7C䉃���چL�C_���_�J5�U�_�pZ�_�����$�	���8�o��R�@�,8��6��hU�Wn+�T�W�J��0�[�tɵ�Fԧ�>H��!�(^� t�7d�@ �(B]��A]J�^����O\����w���`E��d�\��pN,aN$���M�{R|���Q��[	BS��f���g2�7Qj�IǝfZҔ��� Q�D׋Az�)"���:EC���E�̬��m=�8{��Kc���hg獑�6�꥚�A]	D��3���X����@������88�m�J�A��!�����%��~�1���R�y ��)"��l\l��
�f��g�b[l��mZ�[�)�o1,�Ծ��/�k�83?h������д�Т��+���X��#�g�d�&Ф4'�w������J�H�5)˹�&�����:�B#�n1D��G���r8���i��)� �=���>^	��e����  �0�ԟ����L.�Iq�%ʡ�[����6.ǣ�~6��Nm'+�*	ß��;�
���:��9Kڌ���)<����3��u]�v�କ��'l�%�_t��H�}.�)�Ю⹅�8C���8X񒟎�u�w^��mf��]R�e�ӉB�/��r/�$��.f�l����1L�ic�2�P����
��t�T�er�IrE>:�RT=�eՓvc"��?�Դ���Y���F��F�3>�}|�&2��,�PنiR5(|X��Ixtv��0���mJ?������w�[�q�60}�XI����n�ަl%�<��s�?
 ט"��|v�06�g�B��l� ������i� �Ɋ�#����wk��=�dh|)&���*o �e���Aǐ��M��MY=|�0���>O�L��4�+�b�bu�ew�a�7+p�=��;Zy\Im��,��G�4;AkNO^�fSb�[�ߺ�p��I��^T�Jn|%}\@9igڜp�����֫g�~��Z�Np@�ui�jA'lv��-��s���2�,������)1��h[��5f=Ő��j{��joψ�������hl]������˄�����WwLSk�ԝ�v�x�K��n;}�Y�8>?�h�ȫ�^ ��������6��az��(���&���S�S7��g�Ğe�%O'�3����PEA��m35ĩAR�����{
�T���x�'�@���cSt���sZ��3�@��V��N���kK����ӆ���Z�<Nq|2�N��6����z�� ���	$���S��OW������Rl^]��{�3M�w@:	�y!G�N��5<��Dn�Wr<�U���Ax�Qd$��0�ڰ�P�Ʒ<���{���������1�b��&6Ʌ2��6��v���P �z�ʷ���ui���	 J8��w�э`:�e4���S�]�,Z�Y��#�</���Gh?"o�(Ca�v<G���Q8�C@���@�}GAw6��un{ސ�kCxsH�P~���_��I�.P1��*;,Ӡ����ZB��1R G1j\ٔ`�}ԁ� �����m�Ȍ�;{l����ߵ��y:a=4��FO�Z�J������FrLE$�/C<(9E/�t`>2N�Sn3����6/Ja�N�λ�@����y��r*ZkrN,PH�0b��ĽUKM�j�{�fo�����*F�x)�w�m!
����X���r�p#�@�
�&:B�/��s�ZGP�.N��r�X`�����~7j���-)�\1&@4��I��mE��3������
�����wq	w󒞮�5��)�1Դ���]w����N���!�t�5$˄� ����Q����ˀ�x����E�N�r�*)��o����q�L}�p�p
@�����7�eO�� LC!�48�`�< �N�!�Ȯk��ϫp��������Ք׌�r����bb���0dlZ4㠄����r:l�^ Ud��u����c�Jb3K�G�r��Oߠ���uw&��60�y�J"�B&8����\��ү�g�,ݜ,}s=�A�ͪ�w	n�&`�0@9l��g���\J�5�>���Į^���z;#K9�W��H�^$N��DEV6R���D���&#�@<�����ڣG�	�e�1kn�b�_�D%��F+L��q����X�x<��?-�7v$�ί��vX�qS>}�|����?��T�e���~Au:�pХ�a%�现��s�XǠ�k�q_y����q�J���$����\��u+P��u�x��b�U_�?<�ͷ��P(bmg��k��E�蕺t�g�{)o&���7<�W&䴑��a������a�@�q�5�Tl=���������6�e%�+1��w�;�Fn�$�'��e���IZO(��2�q�W�d+&�h�A�R]��:�Ll��w��r��t��8[x��a�O4�HEK�`�D�HV�Dd��Ü#���CDgx�-�R[Y�ҫT�͉��/�uC�d}�Y�{��v�:��_=����»Ʀ9}����Y�x��Wn�H>�`�2�V��k�~|���$��W<�3>����Rm|�Ia�}�f����09������Ry��!N����n;�� ���%���0��#��5@��:!l8�}*���մ�$����Zi8L�Jx�|�XR�="�����^V�J$����Ǚ��!'Q�Dћ��2&�^V��3E��P�^ut0����w���&�ꟳ���o����7�{���6�v�����ܾ�Z�IJ�`ܷ˓KK�㷝���P�-��������/V"�=�<>m�n�|R��%���ڦˍ������[���8�~�~,�(�x�����\�y������}��6��h�"r�F�h����լ�[�	��AK"zB	7��_���]��x.v��q_H%�����Ve�>,�%�/ ��O^�2��699	'kk�gP�,���_���낿��{��O��է��Wk�X�~*Qw`�n(���xٝ�(�`=��_�<^�)��+?
铈v��Jz6i��[�H���v���Nq4�ޝ�X@��;*��M��Q-z�޺,���Eo���d�?�$Iſ`bd{�Y���'��g`�]	���,pӠުVz+>ش�gv<r_�(к�r����H�c��1/M��&��kc1z����lI��d��$���t�~	�M�r��ƣ����T~��6�L�}�(>��q;+~Y������-&`�k9Z�;�Jjn��r�k-I!����7a��;��`�q��gV�^��		�~ �W%}��7s�\�^�4"^�P!Xp�ŉS֧`a�)���q�.1!$]��b*D��C:�~k���EU�h�&�8��m�������K>��s��'DQ�m����0/W���|�^�(T���B(�����)����_��"4�����}|ȣw��HWb�u��b�%Pgљ�Tj�m0��������)݃]_�5��'x�Q���P��J��J����B��ܽ�fo>Ҷy3�ԮQSE�t��"�<�|�J-���n��M-�ih�a�H��-�~o�Q��א�wW���Y�l��2v�)����Y�ˢ�a[�������A��[��v����8��>����~�A2k*���Ro뙄��ڝ�^�X~���t����f����gn��@�����[sР	�?0_:��}�?�s���r���O@�>4�����{<[�ܵ,��581�8�<|����� ���ʎ�B���0Y�;�!��S3C{o���[SFʌ5�6�d$�����om-o6�lX(�Ѝ��|��L�����χ�~įZ<�[s�����;n�F���Ӷq� ����:�m����B�T�: ��<B���+�͍YW�  ����\��5P ͧ|1A8��+���QE���ߋ����P��+	�e�8��oW �b��%��!�V�����j�*-�Z���*�c�N0X@{u���-�R��M��.�}-���V��z��`����a>n[f�~ޡF7�e�i{�a�h�2�����B�N�Е���5����c���y7;��q�9��Ԃ�G�7!\O�
:O*yZ���<��Q
�r���a�d�h1׍�Df�d�V�g�Lo�_s������_��,g�HY�ϒ3�z�:SBxʩ���X1ئl>QϮ'�|��oX�̥>����iW*�K�P8���f�Mz�/+;�/��#)����]7ʥ��D7�9+�f�9x���m_Θ.K���_ٯ�΂����y~�w7���犞�YV�[�9i6���`׍�#�O�wqQ���s�up��[^G�9�	�;�"g�5�6��4@�=D��6�P��j�!�����t@����}�A�\�\�*����Gw�R�O��Y�s���S��hau�&P-6�E�jOog�c����-B��C�(bu���è ��;��{l�i��P]����__P�v���_�nctr�6�OI�����'a�M8}ڽ��y��-�$L&�ڜ����Y����.��X3;�p��Do��o{*v���!��)%�>�;n��ӂX�%Q���;<��H{��T����=�a.ǒ��|H"���:��ݻ.?J��2��}E����f�AS�
����{I�OK�2�=�wOZ��֮Mul���:xk����z{v,]r鞠�4<��0���&�Ojaiσw�z��XG��T��
9��J�ڹ�9Y�xQ�ǯ_n��k���3z�;V8�1S1$��c?΀������XY���DT�2_���\E��aw%-|y�((���9V`s7���i>�����	k�ZB�ʶ��n��J��E��J�b+�ʺX�2*��'�h�{�X��.Hfbb�&1|2��J�Z�C���qǐ,�Һ�(Y�������ֻ��۪]م����5"y^P��ܰc��l�L�<#ʨt`�3��?Q{�y���/C�m���.$�%o���fW��1�L��P+���W����߼�����pz��9��	;?�k}<dٮ�y�{!0��e6�d�M��Yxv���&�Ѝ֧?�bA8���ξ'%�o"j�����h��Z>�������"Yd�uɤ����9#v��q�`�K�������ܝh`��������P1%�o�9���dd�r�������U���>wMTD�h7�${u����F�K�Ŝ��#�No��I��5y��n��Lϟo�>�T�sd1��~���̃�9���)�wWhsP��fJ��π��\��ؖ�)p�h�>��*إ팲�ٟX���X9��10&KOÑ��u�;�./�E������������Z�O�Yʵv����R���{ۆc�k󢹶"��CNB	3 �m.���/�%FeW����_���lzk�� ��ɷ���ѿ\z�Z�z����ZC!�y�� 
�}>S�;0cg��,�%��������x�f��ȉk ��>�o"�(S�&�@��>���΀���}k8�
�D9]�G�_/�`S���������~a�)^!��iq�.,���vBn6�32���1^J^[?���دqq����0<�t�σ]$M������ 0%��B��'�g�4��X�r����Qi�\z:�3��>�:S�rf<�B*q�ء���	��
rog��x��4{���	�;^�@rھ��k���[QG�,g�>����"�J��ij/7WH�]G�D����5?�K���i�x
sz�d��!��I\ps:��\�67����be�͍�.��L��b��%q�g�^�����ޤ
Ck5q���o��">@=Aɭ����e�1�Ř��3��ԉ2�����B���azJ����/�o�gh?-_	���=�$BI���.�����v�~_���3��\���Ə1>6��o7)d�a�����_��� +������x+�?V�/N��}Wl�����9�'J[˞jM��U]���j�j&l�?��ߦ��$?˳y�IM�l��A������#3�4"�%�V�Ь���
�}�ߧ�]O?��H�pnI<�ы�e�����?���U���#�}���r��v�e_'Q�;�#1Э����+�Am�o>�/����O&ڐ#�$E�C�����ݔ�O�B~:���7]�\JD��q�c�E��gY�\q?�>`�L?unMj��p�RJ&p��H�m��:���6��O.��Lf�ç"��^�,qo�h�L +Q�e�ݨ��,�I�2ɛ�;�C�YXb�0�=����S�8Wµ�Y�r�}��P��= 5��%�%dGv{T��C��J�c�jdn0<OM�Q����Y����w�S�ˈ����	/��}�k�c���g�k������=g �K�^�PKD��u���Jk��n{� 0Y����b��׵e"!�=�z��l�o7�#�!��E2{	�^m�}�J��Gu���ҭ}��V+�4>"� �
2��;�I\�s�����'�v�*z�,�O�1��]C���v7�~?z�.� ؾ���ω	�]?n�{裏˒-��/Zy��PepQ�M�R��\D�Į�^*g��r��7~D<$�H��>��{���I����0���x��'����o���[8W*�92�?*�:.��k�n���������N�f��i�;����F�T�������O<sf���Yϳ��*{YI�$*� ��z�&��O�*g�=�Ki�Zm���ك޿�*��pAK.�@�2<,�~D�s��w�_�G�{������%����;%;��*����@�@᱓��Bu�C���"jB�ʇB�Ǘ�FO�C�ͦ!D��Vo�8�2m��wъ���U���`�z*��#h�>k���4�,��nt���lO���|U�G#�~�`a���xI�r,|L�$Zڛ�G�9���%x�w/�j3&}��2ނ�h�S�yi��:T{���/��C��ĨDil��w�޴P��$��=|��̖=����Zw��7:�>�g0~��\:r�8#,t��hx]d{p|��c{�JX㢅�I�)�8�ȿ��h�w�%w,EY�҂����7D��ɭ����>��k����2�Z%����i5B�V�5p<�K)/��H�r�yuy��{p�|uV���}��r����)��[kD�/&������`�(���ThWDg�Q�!5���ϗ^�.Ds"ZГ	s5s���|��!y.�֩��a�`$����׍�T�ter��p�@�Q4�A`Fϋ9������y�f�h�Q'��(b�>��ĵNl n�G֚S�
�I��4�\L3�-S��O���f��lS賴|��5z�oL��ڹ��;�'�b P��
<�WK;�B�K� ��������Q�U%��Ǽ���,jz�M����+ <P��`1~*z3���~I;*�����,�3\��"׷(�t��1O�G[509A��]A(^	3�Yi$�d��-�Â��;�]��N@~[8;�W���jX��-�{�NŲ��{����(��?Kb�Y1�Y�ՕOi3�C0��j�o��X�5w��ϟ�O/���B��n��;:��({zY����	��/h��>{�@�a�GS"%�/Y��*����:�%�b�*~���J��џJ?P�;5�,lY�?�j�A:�R�#һY�/?�cW����Ǟ�)[�y�
<6�?��o�5����
�{������H��s��nh3=G�-�F����)���n��;���_��jSʎy�_ȷ  �ΰb>�LU -��M�s�l�"R�ă�;ڥ��/���w}]fXk<!2#p����#�mqδ����E���3�G�ivX�B�;�A9���Z����f��xv��M�T��]H-~�U�kZN�a'��b-�����-�]�������������aț13�xam��G�K�
g�{����c��m�j�-B鄬�����Fs�Q0��h�U�n��wc�!�0��;*]K���E�Nt���g�d't�T�j���'L[�� �ɿ� �2.�ߵ�j�(ǌ<��AZ���������JZ�b��Z���m��=���Yo�#
7��*q;%���y��Ij ����^-w�UO0��,��V���F����Y�m��s�K��yy�D�y~�M��[���T�=!�`��E�Ƕ
����_��;���r���O�ϟ�y�w0Z�Pc�Fh�5�rsh5C�y��j������j�pې�3�HF�0�(��n���Z8����8�����/��0�K�~0��%m;���r��ƶ�ܻ�J��y�C��õ@p(ll�m��z��v�H��-ܙ;���Z��E�:���TL�v�9ò+W��e�G�\�&(߲I>�FI�,�3�i��W��M�� �Fg��k؅�}�u�ZNz7�{IN3:��i�ń������e�(՞
IQ�`�{g��++��x4U�{z�C�M;�u���]�^�7�t4)�T�������FdX��-����Z�aҙ�L�fW ����@�3޳I�%�_ˈ���a'���.��+C{Ѓ��y�a�8V�8�R�1�kU�1�2rAٓ��I4���xSP�uqf���p<��h����:�i���N
K;�z%�t%�ÈKh���m����3&AF=�ύ����|���Z2!<=��w5X���I�-�(���B�u� 
QA}v�y�'�3Ib�8%��:��S�����;��{AGJyY1XE�XG�� �/rn;	l6��MX}��S�Ki!f���=8�t�'d�:[���#�v6ƚ�����\�Q�B'0ʊ�S�*��]��ۭ�!b�E��k5���/;E�u�4hح�7��G�:��<�Y9}k�/���-v�w͸�� ]�Yu�_�G�
	�k�q�Z�^��u��h?}�"�ת�ޛ�����5fmX� k{3!�$��|ܾ�Vk�OL�QÅ�׭�tZ
�v�6�
����EEj��}��?�nt��*m	�}��G�yk�d�ff��`�9�r;�o��2�,�-��ܱ��tF�a�f�`�`��Of�wCP��]?ZU�rD��G*��~,'�D���f��{Z]P� ��@��^ՇpvQ9n �!}��z4Х{'��D���4̸�շ0�26��ܭ�'�6��k$�&�%�]烇��^.�j�cP~�Dշ���]�T}<��'|�����ź��'NK8HU)��ufO�#t ���KpZ:4�p'�I�I�jU��<p觽�&G���LP�d�"��猒�����ߙ9 @�=47V��u��k��%U�Xh���A���"_�h���˙U��N���F��ݴ�;�]de� ����f���F��#�z?3Ge���q.&��8�6�Vbq8
�!�j7v|�ub=������ئ?�>�h������%��w�5F�� ��J�JB��RF|��X�'�����6��_,��Cv� "R0{��.�T�nQw�{��h�}i�򭖞8?Nٽ?[n,�ć�(kDʀ��A��}���Գ�S� �ȕ�&�
�'�������Gnn��u��ă�G|3Ih,��Q$l3K��r:x�O���^�������t�*�eg�_\�I�#fj��?jXO�5����l*T����z֬˶�uo͍�h8-�q�Lbge\V}xt�Ĳ�@͍u��3��ʆ}���	�����_5��?�4�onԠ��;�?�N������T�%����1��2P��)�������]vC0N��PFW����������x��������4:���������!���q����� �dJ�=غ|�s�Q�u�4�d��C�X�2c�p���{m���l)��XI��ˊ %�&��8h3���楣�58QNi\'���������@3�z�]��t8�1��C�Mf�W>���������O�np{��a�Kb�1�,H�QR��kJ�Qإ��(r3I,-U�Y�s�pZ���M��Є4�	b�sr�:�B��Ч+��蒅P���>'�^�����7+)�_++�qU?��z9 ���.�~k8���>3|�ʸ�������5�4���[ٝ�B) u���tge
�b���h\��R �ȫ�wg��x&QӨV8��dN�s]|Nt���l�D���=��g�a��,
w�f����o 3�<n�{� ���M��5����\���=��*И�fv�KO�'��fa�7U�l4��t݅$�)�����bh���WhgH�G@��4V��|/:�H�<A!�҇_l&�'�]
��/|R�����s�M����uy���g��Wy�ȣ)m�v���z3h2)��45�)?Ί'P�h��7D����@}���@� �[f����{56�#ͦWg1~B�I�"��<��E:=p2k9�R��Ѹ�Cnz��f�QU�hT����}G���#��V	|M�2qa$�XJ˝,;U����f�6ۇ�P��M_�&VxqTe�C4��p�����&9�m�~���v�t�g����߼4m ����T�u1=����.��1�V��O0��@Q[h����F�}��_3�0!<[�ǣ�-�'��{S�&uԂ���J�� l�5��U$Ф|�s@x�L RBj7?�u|�z�,���l(@H���T�����07����.Xʄ}UD�U���_+�9�Ä�6�d�2�l�VV����r��#X��ߠr�\��Q#�R0E�fX��gu� 0�������e�>t�d�
�h��?���44m����6�M�D
�QF	���)	�i{��������8�$��?�����M��UGY��B��k)F ��jj"��u���\nI�V]��Ȼ�\�o��Z���3���EkFw��q|��®���{6��T#�E����L�]#��h����.��!�h;��û��*�>��|m�
��j����3}%v4��ӳ:��C�R�P�6�t8�x�;;�>%|��P>v>d(�h��v'��������t�jZ��F���_�6��<��X� ����,x�X6�@}���<�~��!�o���o�y����&��%iQ5f��3I�ͻƫ����L�>�7�(:LA��(�qw��r�/�u+��x����;�>]<������t��D�����uN�p����!u���E
�������������!O�eC��� ��J���$]-����$�W��y��O7��zc�=0��f,�5���D��t>rbZ��Vj#�'��l��@���"�\@E�Cv��2���u;j+<E�9E��fm,ַ�o ��ο��q�6�RY��6$
`Ҧ�	�$�;���t�,�^=��z��O�7^��י����*����L=�oX��]U�P{_P�id�>��o��r*d;*��t/�2[�6�7�ß�.3ᯏ�0�5�����������T�[T�E��n���Qa%R���Y��Uu�Yl�o(��=���*l4�zk
"�Bթ�����������"G촭F~r��{/�S:ܗ�[�lh/Kh��7�[���~͈�aes���(=�v�\ſS��^�Nz��.~:�Rk�q�V���?��E��7��t��~:3͌��i��BQ=c�K�;�jc��P��_������ǌ�a�>m�-��?˳6h�W��������HK���oG����Ǆ�ֿ��(o�t��A�q��ʹ=�6M4�'7�c�O��*�s����̷tk%�X)�d=4�  PT��	����Mzk�F;��?�f�T�p�&��t���x�:�?�9���9����3+��D��f��(��H��(?g�+�
 �򇢄�����w�,�̌.�����<<I!N<���B ����/��C�:�W��S�l��	�-�ߓ�����p�d�(�Y����N�'��$l��lf�V}A	,��ݴȗ��L:d�s{7m���Q�/���L������e���^�|)�0Ш{�,|~�OQ E3���Ϸ�U1��n�{�5��|(��u�FGk6~.�{�v��{0��t�z�Uږ�y�k�Z=f*t���UD0�1'z�J��~�����[�3R�xk����Q
���2�2\�6@!�j�͕�lr>o_�"�v�H��T�9��XO[!�?�������0R���a/T�T��d	:|�vҠ��*���2���s�"�� O	�"T� �r?���^FيT�N���r�9*&�L�,x�s�z�%xi�y�5Y��h��qE_����v����Vae�{�x9���"�#b�{si|�?`���aѲ]Z��'I�N��n6Rz��yk��z�,�C��m�QU��3P?vH����#�X�j��ܽ��F�5�!C��j�d��	=˵�Syot��v����d�Ǻ��w��^:6z� jGֱJ��$tmuR ���Y���%6�?UO0K4��JGHB�1s[#��O�Jln���~w�3��?i8��[Q���!� y�u��z���/.�"���&9X���Շ�{砏c�����V_s8�5S�o$���FhP�/���Xŏg�����4�P�6����'"�{��_��m:��k�7��s$�D	�����%�iO����by�/��=���>��|	�D�^9�we��w>�fD�n|�X��N����Q\�$�%r��/h�d�c*2! +EB�<;<�>й���Ul�ނOw��} �.��n�y�FС��#���H��/ן�C!I�3��w߶���g6lG�(�~�#T`�ع�Ŕ��L�+��Z��K�4���� ��m��5?��( ������t�Y̮ƾ�����^�Qʘ��l��l��I�J��;�	��k��F��!+h�	b=�����*	�2}U<������Q�G��-g�����2P ��{>���pz� ;ԯ����澍�����P���Pca4Q&/����X�m���
�<K�NҜ!F�S:d�����mģu67�	xS'���l�Fe[1��O-��ՑZztk���h�L8˘l[�(�7{�p_-�}yZ�� Ľ s ��c��{<�k�9�J��e�����{q��.�;�0�s�{������� ��9uy�:�?e�=�/�������}\���
��?C��������&����������+p�&$.zi�Ysu���EW^ns � �h�.����%���s����be}!��-�~���c Yl��p�
�xܐ��d#����In9a?|s���SFR�|BM���_gW3�T��Q��/�4D��#8�FXk���]5Jţ"�������L�<��Y�N�����+C������Hõ{��c��"Ȉ��Rg#��ǝc=�h Q�3���批D2�^�e}Λ�s���E��P�O��J�z�E���U�.ms�2�����& (,�.�Z6j�)��㺋3�
^��H0��䣭��������.@׶��!	�zN��1�W�W1���C�u{�g�op�SdT�ʾ�l_R愯ow���4㰦[l(���j�e���%n���p��F���E���U�����@�:�+��ʰ�0(��� ,!�L�|�Y�&)7[
z��{�W��y�AT#r�4Z�[�(���٧�����h�E�c��.�^�ʙ:}��H�s{-�C�.���9t�-�?Gd�m=iJ��\��J����a��a�����%@��n��k��R3q�/&�V
j	�����#͌�d�I�	�\��	����Pz8��=�l�7�'�� ���5aE�ކI�\]�@�"J`l֟L�*�O,�t�(� 7ԍ��'��g 6N���5(����G���!q���[�C5�� [&���4{�����C��Q�h@�;������cr%�y���QЛ�`a�p�X�@�Ǜɝ
U�镙���5��q�F���˵#w�^��Mbg��Nf��n��#N|_�8��3���?dՕ;H���o��;��S���N����I�!S#aB���"���G�׏������,�&IW�wP���|��&U�a}}y�ߠԉ|�P������ ��������.3c�=��(���8�Z��O�o�3\ʺiD�b�W��PĊ �c|?9��������/�e�����8u�
G�yB'�Տ��)�S,���.(c?�M�Z�p ������gݣK��i�B�Oi�!��\>.�8�0��K���RZ ?23���~`)ݱ���;�LB��:�10kt�g�s���|�9��b���������oQ��	Ǉ�/ �6��8�^��n^���ᗖ����GJ���C��D3���ԁX�s��������ו]��	��;9{{}��i���2k9�A�ڹ�Ŷ��:�[_�)�S����3d^MvѮ�46���B�G=���/�e�Ԙ���tcc����j.~��	}x��#A:��d���k@���>ʐ66Ճ�'x�!V�N!폶_�^�3�������:T�m�;Z>�x�����F�u].g����x5f?1H�pN�+t,�JJC��ĕ����/�Fl���=`���㱽eo��UN�����8}��ik^J6��F��
g����m�;��=�?Ȟg�%�:������;_:�՚t���Ո��)E?B�P�K��ȓ|}'�*�$����㾕���i]%m��2��5���b�����O���c��ʯ.��c5�$q�F��Lx����*��[,����[fT4�����$��߽s:m+�bJ�.I,W"!������ŉ�W0� <�������BHRÑE��(+��f>�1��q=��O�ɺ�2N��*_�v�\с�)��ah���+�a�&� �K�U���9Ga�)W�\�?ƫZ;S�7�?9�y�c��#ַ��F� I��-���Gj � B��qaw��@�0"���{���I?�NX�g1�$I\���E��Qz��1�\����
%'��1T.]�o�G�7g�s� �X�Mw%�y.h.B�I����LT��v�����������%�ķ�W?�w�^�9K,��S<�pۺ]���'|��x�� /S`��8������O�U��f�q����� �`�%�>c"a(K��ڱ�"0cuRS��8���4u�.�$��[���q�z��|o�2��C��D\�����o����sd�%yR����6.�z�Yyp��s�?:Px�oQ��O�۽<w'= �B*��,�˟�]�/J*��oP���8�����&�1�Wj����h#��.FB�7W 7�P����=4�'!W.��M)s�^����F�t�i��S�27�|���?��?P�޼��Ժ �J��q�u��D|PN=u�s���'�e�zo��@�N'���$�qO�8Q�V0��Hx���Ga�ߺ~Z.{ﰹ�X`'�"�}��B	n�Tc�j�ۺ�C��ύ���_8�b�{� A,�v�d{�}�B�u$����P�A����i��N3\o��7�aZr�4��;�)ʇ�T�e����
�}�S5��	oG����;���s���M��{N� �����8�,&�c�1��2������̑��-��-�B5Q|�1�F$M{½��qc���~ى�1�&���� ê1(�i�I�׽�_9��锿1�籨5�w0S���xxܾ?��������:��E�	e���wa�a6�������i[6�1t��I�Lx����K�t���-��=�w �&�G3�<��ё�K$��:�]@-BAj��u=���PQV]o�Ã	�^� �@	2�WK�Kɬ�Q؄�p'�@Y�|ٲ�A� 8F����G�b��6��?L۹/�c<Q"|5���ֳ���z���� +i���jْ}ȓ���Qkf����o�q.r�ZrV�!�����b����
m4�̯A�e����o� ���}��+��#��]8ȏ�5���lw�7)�@c�
Mb/�B 3��1�1���R����7]|z�9V�0��j���z5}���0 D�� 
zgQ�P31���Lj�K6����0������R;�F���W�V�j,�����Q'��}��W��c�����K� I���'H�ʕ�Y��|�	`�EEu�8�`q�G�`2�O�N���NL�1��B�A�<;�6v"�R/�X��P���W�Hh�|���A���d�p�#g�ѕ
�����*@
3މ���t�(�� �K}����5�xPN�)'R�8Dc$�c�R�W�|�4Γ&S����>������c�XU�o�w���?�˚��ߡ��2�[�������u��@w�I���� �1�C9j��%g��ww`=��Eki����nm}�պX����k��נJ<�/Xzg,0A���RQ�pVUH�F$�K�74��\�.�� ͷp\��5���p�����e�b�0�%5�˕��������0��E��9*d6}��U��
*�Q�a�A�RAML�ef6����k)�t|�f$�p��g/�N�i��洝�h#�y"ѳ�-��'��g-x6��X�L/�5r�?9v�+9���8����&ۛ�L���-����2P�s���D��c����mŗ�d���ȇ��2�y��mG���,�gD��xPF/�x�=ypFF|6��y��$�s$L�����BF0_XR����F�y�<��?�&~�%��7j]Q�4�oW�k~�RZV�E��G����[~L�ɂ��Q꤮b�n�pf'R(���w��H�z�����p
���z�#6y����b�~�Z�Ņ�#�e6A���z�ŵk&|�!���"�2������B@��'"B��qh��	ٸ}?`�Ó�hB�Z�GF3�п���o���*D�:��Jnp�ҽc4[Ž�L�,G��ӧq\H���h%|�|�T㞴,�{�T=�1.-����o5gL�Vr�v6��c�p7���!��nNhw?��zE���$���e;m7��W(�uG z���'��}�H��䮥�X�w2��v��2��1���W�����3\eVP�n^�̓D��6�T�Lx�7��y[�FQlDq	K�I��m�@�,o��r�ց\V���|�A�lk���ύ�8']�sǑ7|�?��mx���Q�.������������Ο__�3��0Y&d��!�wN%/�i"�)��3C��u�C���.�t��$^5�S��^���o��i������+Kl���n��ay٧�<�9�U�1�����i��uȢR�A.���X}�Jܧ
q�����&ja�\م��	��j7��t%?M"�h�RZ�
�r3N0:^}���Xt0LxL&�3�F(�g+jE�2�s��I�N��Dߨ3�d�
Z6��VnR9/��'���"?-s�]��ݺm&;T��&ZV�k3Q�{Z��cq5���D���W^�4U]�y^��@!2踶`Qz�����'՜��]ƙy�����C�;��?g���¸(^���'�i�&�1	�#ʵ0=�l6>l4˖
�i�ؐ�S7�v�_s��7|J�)�
�RY\TŰ�'�DK,rN���(��4.�8��'M83�0r(C�uB(��r����fXep%5Hd1�3+r@�>�� ��?�j��?)���'O6��|ص`�_��01�9>�w�����5���><�Qv��q�C�|�P�06YM\oR;J��+�����/���#��tD��v��Cz�,{���Z�L��i�m���h���sE~|\%��T%_�����o.��M<�>g@>�k�QVr�b!��ZR��T̾i{�$�G�G���/�uX'6�[?d���]�<~�}E[��0�پХ�/�9'�c'����7V�֙��.>�ʥ�ER�-@�=���������+Έ�c@��(U��̊�v�#'d��U�'.�pT/�\KY+L]Z�j���b������hIed�ܿ_4��� ���FI������5�7���Vu�:��*�3}�d��/#�}_A��8��}���
�и1����e�ФjN�e��olA�	��p��}}'Ld��Uڬr��"u!.�B���*n�NN[�4���{�x�F	�j��0�(�:|\eK"R��2#�5���MbxV����g����إ�r���M���l�����Q\w�$��R�\cZ�������|���ʚ��y���pQUæ(Y�!��������S#���3�oE�T*-k)N�ΏV�#��}�?:�W��w�@�kyZi��}܉��>Ts��&�c5�������T jΰ`ȿ򭵣�{�!��.w��n�ɫK3/��a���mlTEX<�3�V?�ų��o^'�!/�з�����+�N�o��A1��Mu{w�$%��f�\3Z_�*�Y:ОY�[�Tpp/��s3�t#l��Q�thߪ�	��c����U`�C�W��T���J�O�fp���w?1�tDS���4�r��W ���D8:��q��@S0�mC,A��س%�1R�=����w�g�;�h����5db�N�cU�/�?]�~AS�t8�f�V�ĥ�@*><�]#"~T���0�;��|��hn�J4�W�6C�Pvt�K>K�Θ5�����E���KU���{[��� ��G`��_����7�(Z"S8�*ݡ�k9-��uD
[�� ��"m?�p{�t��^ ��T�����*7O=ѮK�6���*.Һ6Ц�p��N�?!��-��U8�3��>_)����1�;k��3&/�M���Ir[��O�p�΍2+��6��a�X���7v�5�V� ��!yx��'�kc�w��n����L�Bޒ�S�O]Fjb zpμ@�C�c�)�FF1m2�]�oq���="�>
��|�d��(Y)|9��F��Q�.�4i�Js��]²���.�̅�#;>#U]p\�}�b��izd9Ê�ą��n8�G����~��=Q��,W[ꈈEr��/�x��7�-I�c~aGBܬ��@�X�1'T}?���u��K����7���Ŏa�^w'�^����YЋ���T@����ۧ
弯��Y�/�A ��F_���mh��4�Q�˒F�-�t;�|L�<���!P{�'j(P���b!� a���/k0�� Y14��bhe��]��/F���P0��Z�3Z�?��yLx����ckSw��H����Ǔ� qW
)�R�nS���h������s�8��+�e
��i�~�NRiY'	�=E�z��_�H�_J���u3\�~+����a�N3x0���z�w�)9�GN=~��j�kk!3'G�f4[�˟��p��ɠ�߀��^KfČL�񢵷��da^�X`y �� ���Q��y����c��eX�_��g�	�%� |������k�k�)��x6�Ƚ��*U{ܿ�쓑��V��%��r�7u˟+P�,66�_�kR|��ʸh��oħbI���#J2�5��C�+�̿��v2Ė����G{tt �n-3r1U���"���_OV��[g'{��7��b�)ĩ��mĐyG��x�in���7;�U�d9e��-c���Ö	c�wҿ�V�]�_R$�v|���Q���+'8%[��n>C��y
�k�{���5�<�� N�檫�~637�M�?�8=�+��:?�2��.mn�Ww�q���ml��0a�#�h���"rmv�=��s�NO�8���g��0x��5�%崭�6�3K���'w���ͯ�����s �g_�e��M��D_]�ƅ&Pӗ�����
�~��s�T(�y���BX����m�/o�]�Z�0�ȏ��C�{G�EY�<�4��FY-�*L���A�����}��2���#�`���nyq��v���
�"p�����ٯ������M0��,>��=��!�s�*7�k�ZY[-'F[s��9:{�:0C���lZ�A��䑆�^�"X�3�J���ԣL�ĭW�V�+Љ�l�had�Ɉ�9dxt=���W���dEa����9bFR���jM�H��4���ޖ9X����'��a������
�e�����[m���~6��4׉��V��z�%C����*�܄<�J��̀�p�8�y�-����m��Ķ	��@�t�	�[蹠.'���B�GK���f�+\���E�MUa�}�V���Rdk
��WTC�.��V9����*�Vf�v��9��7"c�-�y+��aA}kÎ����6_���ʕ��{�X�׸���~��y��L��F����P#�C�`��p��	Z�)9��xk�-2�G��r�o�M�m�k x�*r��=�i(o�"�;L6ف����D�H�����^��"��(O�?��!�ʪ��� | e���#F�i٢�*�|ޘ �7_�o�ݔ{oZ���9����{�qH\�(�>�!y%���hG{�w����l*������X�?N��.��ς<[���[�1c^~i�F�V�y��u:�@�b]�.L�A�IFx�u�s�����	+�Bi!�O6�\��?��� �g�⫰�ckk�~R<���&����K>�C�@Y6��)��>�ݖPu��zE�pf�3��}q6�S����0� �ӷ�t
Xb��,)�H�o*K�n�t%�{��
[��ū�˕jo�a�pT Zh}���M���qǹ��V���5��� K��3�Y~Ќ[΅h�1�fu]E�z�
�>��$)�M��[��Y�����v�(�0,��!*I~�E��{���$*����;s�
�1�=������Bp0#����ɁL�v��S��q�4%%�T�~;�D#E��j��"H�·�۞O�-
K�ad�ٕ��}@%����f�$�zk�����5�/��7#G}i�]ƣz[���D`M����]�E����q��V�i>��	����HÑ���Y@�F��D{;�8A��Ө�����!μ}\����I��%l[L.�R"s?� ���%K?�S���V����G��/�	b����"��}�9���5;��$��Ra��YI6��#���:P��ɮp�^��II�A�@(�y�y�P��V%�阢ITpc�
U������&��]��B{g��#�S����f���``���M��[��Ӏۆ�O��k��$/�-�:e��u%�%�D�{����jQ��~)6�p,,j���ON��:!K��54)6#��,{��	���b���#��]�(��t�B���Dc�o�H��d�?+�Eڊ?�U���lS
�,�H�y�+���CgpDʎ�L����,��K�x�.,�N)��߻ [��j1�٭��?� �0�=�%RC���a�ɊXP۷��3C���r$��H�*����Z qmo�ʚL�2eϽ�)�<Ľ.�N��.H�b),��1� ���l�-�J�RP�3k�D�QO���"�E���È-C������A�>nK�L�)��}TD��K�0��%��!�|����MR|�d2�u%��Z���#V����
���Sh����'��t�-�6c�0��B*{	K,;�����k�8BMQ֖����4p��� ��H�'���Bab=-Y=L#�bsN����[D�Z�>��P �`b+��󚈣o��=��d����r���֘{�ۆ�Cc\��[Ms	֯�E���.G�?v�u�y�$v��-I�z7V��/�]����h"�"��7�p,�)�R�^t?�3���U�\Kd5o1;���G�����ωGb%�e��Y���Kf���^��m���,���)����T~/@�ĳ�^�|֤g�x�rO�|���4�	��jq���w�卹��%l�l,a���*�>�`s���JN�>P��T��F:�F9���kǊ̳q�B�x�h�f{��.{ܾ���rð��Bc�4ܱV�5�:Ӕ�A��Pc� ��/��`{��IW����rډ�2�P�y�ǉ�ri0;��1 t<,�C�P��/N�l�J۟o�T��q���)y��$*����=��c������$�4I%9�Cav2�� L���պ�/Q�>�3,��R�m�5̓��&E]�΁����Y롢>�����l߰�D�����D�P��:E@%(�ʳϻ,�F/�=� �GrP4��[zCv�K�\�4�RE��B8��B}�N�L��+;��շ�zG��̛�_)��]2
������켑q�E؃G�|�c�pk���_��,MY��|�]���B��F�*�����8*m�~���EA�	|���:J��@sþ 2T-���L�r{љf�%�8�h`IrAރ�TI`�"̚�ћT��p�'�T��##�_� '�A�"�����Ϫ�w� ^@/#l(	x���$�kcyLiLp�}�*�Z������):����H*�����q}��M�4�ʤ�oZ�ڒ00����ơ]�!���K�b��B_Q`i�+Qp�Jq�[���mb�<��|�F��AkFS�@�����S#�����jM����hO ,�?H��8E ��p]�(�k���.��Jl��_
��E%@f 1%�M�O#��T�d1�d��Zp��o4d��q���a���g�h�q�?�	�y{mɫͱ�����'�
7��#��بc[��[-�D����Z.S� �]�u���ԥ�d��<��hk���zs�X�:���s�H��m�����z��_�M���M�~}8���?(sk;�8�4�;%*N��E�rT����0�Z�$�>QU(�[��=�ܖ���g���}s���qI�^���JkyH��M�^2G�ȸ���0@�s�<Ґ�����BIBQ�>e�x�\�4fmd����BS��aX���t��e�N�w��W�oľA-��9��.�wX$���a�@}�S�0���d�o���.�����~�f'B?m���hƍeaqI^3�a�N�v��鑎�(`��a��� 4CH�J$���u����7Ɇd+D/S�]�3���"D�����F}~��h�-��t�޺˱�q�jQ�z��H`j��
Z7M��Y�����)"�:	%�&y9�b�dy�WF�-���1��}c�Dw8�&���3�gc�� ����63�h��O�y&�u�����}a?�96��۪�S�ݑ�/��Ei�[�����B���tN����k�<�ѕ�ٽY��0V��D<,�dد�
�5�i��#4�P���r8�>����ɩv��FP�zw�ω�P"�ȋ͠1Ӵ,Pņ��(CO\@IN9	t��k�ĵR�b[wy�z��/�CW+"�9/���Fuq��PS���b�)/�M�7�O(hw  6�4E��n2���-Ž�/7/�NB(9�h�?��=*ldn��L29����@�l�_2!��뇟�CI�L<���ާ�"e¹H��ys�<5 ����V�q�3����\��EѤX�ni�Xc�2�S	�Ohm�1N`X���hR��z*�qP~�x`�C����ǿ�Nj �>�YēK�Ro�4�,�����R����$B�"�c�;6��0��J��u0~�}�Z�{c$��G����*âj����Hw�<4HwK#R� �C���!��-������������w���Z�v@�ގ<�Z�ba;\��2�JK�p��� Gn/����� �F{���[mi�ZE,��8@�����~�"����\���@�Xb�����6���� �3���}�I���c9��h�/��� j�B�C�J:�﶐��2s����D�Q����]4CW ��xc�|f��Y�1��CI�܂���=�i��ω�,��h��nn�LԷ�B�t�����Ĩ?K�6�e+4�~H�1��� ep3�RO'���C!](�(Qt(y����,�D��JJ:����<��}L�
g)��F���N}�����y�c\�ss��c�L�J*s�P?dr�[�D,Y�T<̫���Y*�>C��Y2��ŝ�_�aW�%�:���ۋ%�|�h�.[�Ǟ�L�"yx}�l+�td�	Ry����aVх�?C^ P�Bo�_g�ҙz)����JM*E�r�ܗ��RQ�o��՚	�ȃ%�"����q�h�ѳ�4��0�,P�:�L�Ժ�����ko�
ī8�Q�����~g���L���b�>��@lқf�pj�s����/������s'X�LP'���яƝ� ��_B^[ݝ:JuD�ؒ�pK�@�Uk��P���4���F����$�oK��{E]'��T%yM�cy��h{}B[Cx�F4p���`�yE���8!�ó��ʹ)e��vZ��p�͠�r�Y�8���	��)Jr�G= �@H)�Z��=Z� �:PޖTR�@t6�:�?J-���/���0�������Ibi��E_8uMBl��
>!��3��2��I����f8�\���lB��6�#��g�R�0���S
�'7��ru�r�3l݆8����G�9��f���n�T�gJ�e�7�鲁�����+�TmC�8�q��Z�^�b(��-|����Q��X��tתJA�g��ܜ*��) Z\l:g\����M�tT���VZ@p~�u驺��%ʡ��4d���kC���m���%Cı��Hw/��*8nG�}���i�P�Z��
���&�&�>*�ryDLU#��p��[�@^�%�����O��\.Bj�VMM�-6����r���yj��~oj�E�1��S�$X�m��b$F:v�W���rw��x���Ls��՛�t����%�ƥ�z�#S�6���p�6C���ɒ`Id���jg�ivQ'uuZ��������XCc'�X�����-���:..Y����r�󑗴�<�2 �=v򝠳�N��~畯_���	$��sD�i��=q5rJ*<�K�vw˥QR�)8iq6{��VA�Y"u�/f��R��~kZ{s)l�e��V�
���FP��K(U�C��7�C
����D�GK�b��a�8g�B����:P���|�v��%�U丨��叾�,�n��%���1�6ˁbbY. Y�UT�����ڱy�ꚗ�j�,C7��hE*2�K�p/�d��:�^C�;�P�s\HA��npH̝_�j��t����y���B$Z�0��7��,�[<#�x{Ԝ"�����w���S2E0v�gpvʒp��|��j�M-7�ҍa�F7pu��-'w�򳬌a���a�,\�?Ka`�f�Q��r9.��#G��(���m`��T|!�˺��q\3k�w�6�>u���c:�s�͜���9xB���p��v�G����	ʦ�:�qv6}m�����y�Q�f����M;���41����%5�k�z���8�Bs�b�Id�����r�
vĭD�;�~����I��Ze�R<�_N��]i�T*A���l'�[�F���^�Z��Lы�ۿ@s,�B�$��;���	�lkv]����Oo���9�5�+�/w�S�}�M��C�e4"��
�FlKz����=a�2޲k�v{�stq������k�<�m(c�~,M�i�ٯ���1@�d�y��Z1AAU� �V?WrH8���Ԣ~������1����U_�Oϙܗ��lηN�?�zW�x`Ɍ+޽8x��<���U��Ɖ'hk���W'�s75ظ����䁯��ݘ|øa�� ��;���t(�84x}�-��cd&�8B�n����Ku{�(�&�9-"���Jz:��Gl��<$4���'0����7"�c'��K>S����˫I��%K�{�`x<Q~c~׽)���B��wmΙC��/�#n�[�<�i|��=�$�y���X�PI�v������"M��`��``�*�����Lm����` 1���]z�cҽ<d���[��@�j�����x5����g<J�G��ȥ��~�E2��ڼb�'r�LY�OE�:Y[���S��_�[�m2���h�M��چ�卣ډ$�� )8�v�Qo���t�|n	2[�`�ۧd�*Kk3�+>��΋��ǳ"a���,���ѥ�.��-��#��.�1H�	m<��g+FcÇv����lwjq��\�.�̜�u"�{�J&B2^���K�u"w�Z����R����]��x�G��������	�c�o�i�e�I]	�wѸ�!~D�46kw�&�yr�z_>�.�mEU���+�����?�䄎�/��]�(�o汦�<�C�)ח�?D�܌��a9��Nk��MU�P�.d35�1����j�bn\J�Ĉ�#h� l*L� j箫��X����]��Դ��4y�J���9!R��Wr�����*���keȹ{�J���o;{C�����Sq��Kl��z�Q�sIf��ͦ!��"X>���s���7{�i�m��XIOb�/E/���Ȥ���g��i��ɥ@���t 	;������h`���x!����]�S���v�C�u#��"�_i�M�}<z�_r��$l���L�_V�f��$`�OǾ#I�q6-�>��9�5��H���Ŀ8�K����yyGћ���`������|zg�i�~�����*���S�+�!��v��F|x��Ŧ]d�O0o����/�Z�9�QFK�W���*��5WU.zwr�:���ad
}q��.m�B��G~��@����l�]�'���r��;x��@��u�:	�/�B���	����������G񣰚5^L��+ݬ�s��m�`��D�4�L���0k�aB�;sQ5�1&�Eʜ]?����z�����:Hb��˫��^S��sB���2��>理��h�����0�8Y."�-o�,��>��������2�����-vxo˜��#L���3Q"[A�^s��0[�ݑsH�Pޫ_�q��S��ynNo�X�n�/Ǐ���M��U��N���D���,��Y����;p�Gmn{��K�F^=���U��X,͖qnU�m8:d8�7��A�7S��乒ޓd�pV��	0���2~�]�p��S;���Aa^>��cZ`":$�?d�'�c���Z#�-�ܰ����0ʑ!���^~ ��bŤ������������[3���MΥ��S�[�����*�j��xcG�%�#8*t��@Rā���07�����m�$Y�Os��4�V��W���ҜEw��L�aR�PW�#{�0�g,��ZI>�Q���Z�Ne���X���~O�(�ҍ�g�7�Q�H�g� ��Vҏ5`����ǥ�)C:�ۿ|k�� ��m����4�+zܧd *�Gl?r{]�[��Q���^�ҏ8���m\�} �l���tv8��+�扙.�@Y�u(j�-;>����O?u���9�|�a�Jm�0��0F�(��
�2e��Zƹ���?<�N��I���ugr�Euv�e7����Y�&��2�~V̾`UN��-�����
Ga���e�l~S��k]�S�K�����>/>]Җ	�}6߬�4dsϨ��6L�Ǿ�>���r��U�~ɯk2��>B�vA����-5��W_���,���u�zT��k�����6��	��� ��ʌ��'.$c�y/?F0�v|�=���i���q°ed0Ե|����-�0�Lp~�[�~\��`�=�hQ��{[��ȗ�~8�����!S���]���*9ӌ4�$�B�èV5��O��H����:�M�A�zB�����������+�wANry ����4��wr��4E��76�*x��PD���F ��j-�?������E�@~n�MXWA��g+��
��J�{���o��&xA����~U��+!&�~R��xɊ�Y!�\JNʭw�M&}}=emì�<djy�N-M��Ƥ��y�
��jȍ�'���ɮ׫ڑ��(�Bsy�H��qU���<~k7�|���ģ�����\0�|m%�U?{������l9s}]"м��%E�b!�:W�/5���͜Ρa׎���G�6�A���z�ơN,�������"����="�7��=�+���U���(�X�Q��*M��w���ֹ	[Г]�^ �V��0��5:������ �v��W���XI�)�T�����"y^Ya�a��³����Ǽ-q�ߖ=8����P4�����2<��H4�L�G���܈�w��~)[�k��A ��fw)���Ǚ����;	��O�@p���}&���S�o^Ա?,���gyx�i9��mr�M�����cP��$��$k�����R{� ]��
d�]|y�k�y]��*J����ʱo;b�[t<YPur���jVR��x��o%t��*��u�����(uIZ�9O�,��"Y͙�E
2����b��e[>���^(�щ�2��)֍h��_=�V%����hv�0{�������Sb��^�#�,��b�k�TϷ(ȟ��Y>���Ց�F�����1�l��
=��;o'��<�]�9���QV�?fC��[�#�R�������2���Һ�?�-����;���A�ɽn}
���>j*����6�O�OVX6O=��{wf8�P��=H=���� ��K^�9!��T2�~�f�N�u�2T,��u��r�!�u��e�a�Ur�'F��;�B���/3E"��``o6~�w�8���~���b�>8-���(;�_Z��H�:S\8�!U����Ȁ��*ۓ�@'ʕ���f�Ҙ�&K��G*?w�J�дC(V��-����1b�FCQ�%h�tSQj(�
��o��_��6�y�_�Y"7eZt�jkձ��++ܮ���b|�&j=,j�2s�^����C���<dG�㦕�HX����1��ڔ�K���'n٣Z7\y ���������Q�J�Kl�@c�-�'�íw�>�=��Y�%�W��2�l��YD_0#�W��/_F���+�
1#�_?�{�=jaӽ\���"Q�$���H�dW�?��n;bX����	O=�u:�^�U޷v��$�B+ʲ���=�����������ƼP���Z/�ʋ�U�N��ELR8�fܟ���x�ڟ��\z�u�?0e��YS8p�]��N�]��`M�W��
�h#a�@%m��^���L����}fz���R��O��e�c�4�x�$G�㙲��N�9T�b��B�,�,�x���4P�7��6��f��:�v~j�F廘�"�ҝ���ƛ��c�n�Z`WAJXe�l��a��h�����fb�����-��3��U`��?\�L���<��F褥���!��޽$�NEC��!鳹�2�E�����׃�',�L"L8�K�xV��x��T@��Q���K~*��J`7~�r�!�����|�B�r�j��5o�k���Y�/.�S�Q_������D���M���r��,k���Qg�jq���8N��-6j�	�B?�Λ	���T]\�"��
�R���o%;�j�o����/�W/V&2]�g9Ռ��[y�^�4U?��>E<>�Wk��&ã�	�F_��d���f��!�l� ��SA �@J�3sǉM���k0$�����Z[0W��}��O�A��Θ�v��Z��SϗG�q.�GI�g�j&��:�P�KH�P�דcRO��+�����1i����ܻoP��!�&�j�j��Dx��Xv������w�!������U=m��VtkZ��C �s�ͨ_���U?���VA��[^�d�._5�ˬ�D`XW��Gٚ!���r�+|��B 3��ͼnN �V���,ʟ.ߺiO�EV��J�d�0���v5Pg����(���=��ߐ�%�{�sz���d�K��r?/����}Sw9�N�}��$�e���>����g��s��Z ��-6 ����ѡ�nk??�?A��Uk�$ r�yQe$-\�RM�M}3WKYH���_Y�X�Ω�E�6h�Td��F�s9�W���?��7n�O�aTǥ��#q��]�%b��-�K)'�<"��"��=Ef�P�����_G��ʒ�h�j��
!M�����#�s^��M��X�ć��v����E�eb�ҁU+ʃ����-;	��́�����>�}��6�U8��鐰fߚ����S�?w�@Qe�}�x�l�罢��p>(k%ƅ��L^_jЫ��.C�-O(?�v�C�,�s��uG��Yms�o"s;N3���	��^�8��9Ujm{L�/�}�SL��g���������@8�C�y��x��<z��P��[ȼz�lO�qt�\�����L�ДZ�������2�LR�<�L���mb,������cȋ7�6����%���9m��U���a��)�@2��e�G:�g= ��KF,�+�!uxc�����z
D�F��w��;�~�$��V�r}�@�'��}�����a�%��Licޑ���^$@M���2�ϡ�ˏd
	�y�=��U��u���AQ��p�4��6�p��9d�'��S���_h��o��X96վVd �4�@)z'Q�D�6)����"�%�[z$�eճ�z�7����^ܟڜ�y��i6�JV��<k��7T=�]0Fr�����#H+C�k���
��R� �$�ݘ�]I�Y�K<��(?�s�S��3�gp�Ƽ����",rw�S�Z(�����u�zP)��k���Ĭ�6׺o.(xe&��=οQ�ss˝~���n,D�4>�:p�	�a�~��W?����l��Rۄ�:�Š|9�+���dSy��X�����
���΍�>��W�$PVt�_���6�I���Z�pz���ؤ� ��E��-,�?��&b�u��Z���^
�*����̈́��9l�8����O�o%0"	��k�by��hck�q�4�C��<Nvt�!��(�$<�F�ɰ�#�����U:>����m\�,q���P�46	�h#�&<a��F*i�ʌ�$�"�4���k-���qj�=a@�GU.33��H-?�F�9�Z�O�h��k�+^\�]y�lɨ�£(M��Ǩsd~�ͺ%O\w���D�������1�`5+�F�����Q.F��7"��a�d��yj��KI�!��$���ԏ6������|'W_x��/�($1nt�X���1BY`#Y�h�O��(�W?FB毯�""�:�J�[������N���z>�ʵc
���5��i�j�1�+o�iPb��=�OY<���'�CRǏ?X�����xq�=���-Ѱ�1n�Q�}���/6|VVM��i
]ֺtc�[�� S }�%/o?�C��d�{��Y���G0���e��g"
D�SQ�����agݐ�R����Q*I�ތ�X��^Q^"�*9���}��G�����f�Y��XP�,�hty���-$଎�Z[���,�H(JR����G���&�u��gxo�N|��
��5�ܕ��b�2su!14���_65\���"6�87��a�<o�"� ��u_f��4M����݀�,A���Q��U���(%b̓Q��_W�b��\�0R�������ne����c������x"�� �M�a�n
��Eok��PN��O�����m�b3u!˄�GZV����D9#!��'���Z�X8\H�HK~����������v�Ӓʐ�����":\�臤�=�HO�q%���ߵ�2Ʊ8�#��Tz꺿U+�)I��a'M�{��(��?MW�R��2��=Ɍ�#��P]|P~\��Y�U_s����p?����&�-��֡9�`���:��Y)�� |�G8�w(Qw��n�:k{�a4;���)朞w��j�(%di+�m/�`���oi��lo{�lyUr���tS�k�W�Պ��'7'�anЧ�m"(�F$\L�,��vj��X�W��k{�LU�,ɨ��Ct�����[��Ĝ�q�kZ[���.����*��m��O�©��%���e)���@�X�i��`@3T��h_�����'$��ZB�ّ��o����?�x����0�%z��v)A�pA�Z`��0��i��VY�1_�0z[��%X��x5��\�3��o5*�wx��Ƚ���	a\��c�qs�2�������Nĩ�a�gN5ߎ2�4�G�zo�������V��6{x^�Ώ�F���~^¨d��������>������VݶbN�s�&�����G,_�K���מ+�����L�ٓUP����F�@�3_��\�sW�R�c/��CV*�L"Eޘ��>��g�1Mc�q��x�V���!T�n˜�liO.���*���yWiR��U!���^�+n[�u��Q�2+	�ū�k1�Z������ؽ@{2�V>f�Y�>���f����#���X����ͨ�-Z�1�Uw���[H��X1�����޹��n��n@��C��4�z-9@����Y��͑�f��N3Ld�dn�R��c�cD8%���#�>��:��ia�W��I���[�Y�6
l�j�Rn��)q������JrPq�,�������}ڐ�F]�c�P�XOS�<�s�3&���l�5길@��OL�5�^�6�������k�R^�xFO$&'�a58v��k����He�2��)�u?�=&�/h �\�f�H� ���Ì�$��Ȟ�u���������M!�6�Z�bT4�@q�BU0��]��]e������2��������ʩj
�&�&0����+w� ����R�C����wN��!�7F/)3'��3'��A7l�h�'fM� :4˨\�����~l)�����rԧq�CRZ �I��ȼ�;p`i��-�4	4����Fvٔ촕�6��J�#��Z�`[b��ڶ���#��H��K�6J�I��:�����=�E(�|������¯�r!�-��+���R��8�~�\"�D�a��p���%f���H�u��_:l�*�Z_��䍲���~XJ�C��q׃���b���~�����IW��� �¨0�qDb��⽻����D�@���%��+���h[Mz��>��t�����xL���bS��NF��7�����y6�#b�e�`�̶�u����y�( ��"��'�ibz^�����Qz�eFcu9pX���T��*�̾��e/�~\%��������
�
�VJ�]Y��%�)R|���h�*Y���c,|0=�����{	�CB�r��|��$�G* �n���o\����$f,�����뇆<.#��F��YY��L�,��f�\������Rԋ�ҧ"��j�)i�Akհ��a6R ��D���oKL �Ɗ�f'�ϫ��A��N`STy�v������
?���_�p�h�AD�|9�<�����Rgc�0�ls\l��U���m���  4���O�Ǘ�!�;Mr`@V_V[U�v�$�?��ɠ�tp�2�e���k�z�<l��9Ϧ��ܴA��td�Y��	D&���@�4�"K���XS�2������M���H���9�|����ѭ�;�?����LJ&�CMrY���3�'����y�~�p�����%h��K4W��O��R��;�z�v�e�����`�Sql	�<Ӳ�ߟ8(�̭8=zHyJ�-��\���*U��ɖ�z�څ�.�d������y�����,P�n��c��WR�f4~�u2(�̭��9P]��� ���-t�m�w�MU?�r4��$����v����.�V����WG�K����{`XbZ(��p�C�@g���\!?�+ΗF޻($�~�^#�Bt�o�vr��M����JNEF�Rc�*�?�;����"}j[���c�hh���H#��Y.�>���	�ˬ`��t��ț����d�����"ϓm|�J���R%�ue����V�|j'�t[_�dY����� l�旚*RvQ���P���� U9\ݨD�{v�K�6Kďc���5� �^�������@�D�$���/���w2�����G�g ��Ȯ'2�����g�@� ��*�6�Tn���^�뚣g(�������DX���v�eH�wQ(E����V� b�n��\Ć^м���gƫ�Q��r�ޞD�ݕ��XT���RXѼ"�����Fa��ߢ�M$��yۙ�ի�FE��ew|���a1:\��&L�k�>�ѥo;�(Iy�M4��6T� ��]1���>��YI��
�垈�z~@$Z��W��I��]���iy?�e6�?�h�"�큒��p���?G�v	a�4��XF{�+��9�Hf�sŔ���ǂ#*���;;f&'[�v)ʐ-�ƪM=�zn=�yV��i@V�20F��9xt�PJ��Df��Q� 	{�.����*��S4>�Q��ޝ�h�3;�>d�5]�O�����}��K(4���Eyt�5T���4�����۴)���8:�W�-ޓ��v;������_��d�z�z�&!,#9�&]���iA��T��aw��U�������YJ���F��+S��X!�Q��3��߶X��b�u�����AKq�5�o=��F���B��ч����[��=U��?��E�@i8jm[�,"���*R�O��H=�!Omw����U�_�:'���b,�L���	�\��\b.��Z�ZU�M&�=҄6�7��b����q�Z!XږƵ}Ҟ�N'
 	��oLn�@���� �tΟ��l������c=I�|{M�j)^sӀ�	�:����w-bK@BQ�E����-�m]�5��͕<9r� l�N>=���1�݉��C]Q0D�ř]Q�����+GvU�������Ú� ��8Y�K����G��׍w�<g���2����_�
�_�)��`�׮�n�o}\��@��IR�`M�����+�[Ű.^���Q����x.,��C)aQ��K�K$��������{�(����Q@�>���|�_����@�3�t��V���n�jJ}��٬�����n!yӻ�u=��Zp��3I����U��*��?U�e��S�1 �R����sFny���������倓�Lv
b�&���+���i�G�~��G�zα��vҠ]t����$W�g�_<$�*� ۭn��k�=
����v	�D8�7��b]�M��In�D}�.��C������L&�N�U�d���&}���,-5l��C�Z��'�	\ �@�[zAihmDpC.A�Jؼ�m������R��`���e?�/E}9x[2�:J�Q�h���rT6��D�������~d4���u'j��-a�� �O F�3��7��_ݑ��U�q)F�����uE.�ah��F���{�
��W�4�$lk��$C�F�ev_Xc��~D-E����YHK�|e���Gü$�B9q�W�{[���[��*��НW�w�Sz1�
�۔'�P"�R�Zt��������6k4�c����:�`�ϲ�l�@��('����tZ�~��0�ʻ�BX��s��]��Ti���22^�w�VRy?���"��&Y�;3��Y��Ʈ
L�{���}�6��2����@͇�۱���HB�_Jv>ǃ^�b-t~?ƨ�GP��Q����5�M`RM���**������Y��Tr�K?����	��a�#�V�΄�ͫ�L�~����U �T����ߙ�E�1T���,zw��yv�K�.�����P��ÝC���K��`��s�s�;�'�G�Il)	�����o���&����8U���L��/L�H� '	d���H�I�1���\Jz���C�T<��;�������K8�bU�8 ��7z�#0�B�F��M�xDq��>l9����s^_~��:����͗$ȇ߿)��q�P�V�y�t@�T��&k�?�T����c����������x��oP��i��6�$�^���D���bX���?Ioc2"�Z��/Y��&%7t0:���q�PY�wf���^���헃(QG������o�H6s糖=�^��\rpF�5�P�w�����q9nXe`��pY�r�P��y���4���ʀ>5iz`��"U��h�5��QI�!](�{�_��Ð�Д��׿�P��
���YmNx1�R�lxxG݅_e;e�x���ًT��J���@�d�F�::H���h��L�V�XL�0�ęd��]��I�P��[8Ocs���r\L�d^H�o(�ޛzT���X��5���`!��RS�<�#��I'^_�+�T4Q
��v{H~�����O��(�u8��qL��,7�z_�6�����lx8��,o�z,G!�Pr���]�bF��s����DRө�|ù�c	��|@)�Zw󾽖�&�S�U{a�q{V#)Z������HA��/��oO���qB_9�u%w�%9��x�ft�5}����f�۪����&ƜoZ�P �d��Fv}�O�#?��&6!q�$$]@eN��;/���QG��JP���N��gj��6τ��6@EN��»� �����g���-���4N��_

�L ��o���7s����	*O�`��s ���x<�>:�"�����1�se�`S���ݤ��l���G1Х]�)SF���~z��H���n�ïh�$�hO}@y���>.i�V���M�Z�h&+�</gF�dJkЛaR�l����	3�pI�2>r�~�z��!��2	�+_�f�^d,̞qG�[X��}�nQ|J�6����b,ܞAOtsx0�/y��,E�����GH9�����.������ʘQ���G���7x�-�j�Y�U`(L��3�v�<�xK��,
M�	���a0/��-Z_����w�Y�&m5��(���4�9�Rv��g�o�ovL`��������cz���x��r{�̀$��7��~�L1�V�S�����o ��%���B���,����	A�Е�N��6�?�������ǭ���r��i{���P�Qy�Μ$l�	�����Wbc~7��k@X���)H�N��LM�'R�F�Lp\�� ����<W6Q��p�l?Ѝ�`����'�@=A�j 3�!�4���z"s�D9AB���%9)٠-�fܿ�jg����3pSG���U�i��F3����JoUU���=J���F����/aX�;gW�BiVq]^ѵ�_[��m���P���il�N����$6^<Ѐ�ⷧ��>��jh�$ �
�>���˙&rYQL�~�Sk������!O�R�_�/��� ����f+G�Z��p�sW� ��lސa�v'2�>5`X"4
"3���H{/u��j��& _����Is։�@R����٢�J�a[i� �(��^��� �����g����w�5�'�g
�F��R�p��K	���N!��`�'�y�7�yAt3�?�~z�*�����,����o��9�+n�O��i݊�P�1��c��К�7,iԬX����%�!@�}�lZ�\J�����~��|V�q�މK��䝷�"�[���.X�Z6F.��a��?����q��&�(��҈8���')r膤�|���_�Q~KX��N�$.}2Y1:V��Մ�uO��0 *,�H��/��
�w,j��P�lIYcT|E"6�U������`�03!b���jI��^��L�ށ�$���#���-È���ɟO�ޑ�&��{�CK/v�,a����~w\�,�
߶���o7�e���ӓ0.�Q�bu��,�%Z���y%��2n�~ZBB*�� *{,&�����86II(D��k��e.$��g0I�`rZ�cQ�H0���Ad��5_8����P�k�Ԃ'������!ڋbЏ6!	~�ڽY��u��<�)D��R�fU[&'	9+"(���G��q"+G� �c�9F3�F�@8��4�����s&u����@h�L��{�|�}���e�]V�U�+7��<��2#ʔ��U@fh���ud�W��6hIe��{���Q�ŧ[A�逻��(֌�����<$�Qf��GЖ����[��b:��*�0�p�����w��#���.�W�b�1�a("�M�W5��E:�.v��`%�$���I�5����[`*Q��l �q�ڍ�:�v�T����p�ڣ���p^�0U��2Q?5B��-��n� �|rB��g�$#����{�?)�>?�$��� !OBW��a4�yR�yV��B��u���"*��-W6�ݞ�Dz��v��7v�#4��y�1 �fm�o{������_�1��E*^[�o�r�ѽ������S@��F��v���3��8o`<���Q���W��؜<Dh~���U��������<��{y���)��sGD�S��T51۪5u�D���Ƴ�>r����Q���F���(&�lF����'�+�Y����E���`��u�.�֚���D��b��x\^���+�{��%s�/�<��Eid_��;R7L�	sR&~�^l6ڨ	,��X��ۛ��WR�p֔����U�A��oI��IU�޾�U�%��	�fw�q�j�+���p�[���Kº֚-
�"*�6���me��蛙�*�I
D�S�/�_ ���,�!����7���XD��G,��>����� `��gW�4	t���x��Ǎ����@H����!�Ϡ�Y� 3�_�@Lp�gw��GR2PM"��R烬E��
���b� �ɽg�9m2u�<�%�q�� ��F��? c҅D�ꙶ��$v�����8 �i��$���b	�\)"�C�Z�X���Bs�]<m��2�I�%�k"��/.��� �f{���z�1i���.Sp.}��
�mD��<��) ����Pf��X]��i�`
�� ���^�P��~�����ML��n�����K[�(W��R:��YƚnÛ�e �V8ߎ�i�4�͢�Sh^��T��_!*Gi7�i�Ξ"B����}�r��K����/���K�*������Q�K��o3��3���<av�_\qq��w
��O�@�风ә��a���Md ���[q�&����ʹ���Q/Ox�Kls��gr䲾��L����j-�q��C��9�����ᄺ����m���;�(Z=�4��iH�ג61@�?��| �
q3S�u���}[?����.��x1t?v�gj�V���n��ɒ|?��a�ط�m�4c�TEvr蜋G9�ng�<A�^��Z@�qS��^��T�)��w-XSzd�,?z¹\��i(,I-[�ȣ��@g��ﾲ$���06��#��Qlx���:��/믫�F�ާ����8b{�a���,_��u�il�����n6]8Y�t��E�Ѹ�Q����IVD�'*g��8�(%�(7�N!2M/�R��C��R�+����i�z�����oˊ˝Jf�����p̽И�c-C�S3�
����2��ܫ�E�Q'x#�>�D��g�j�{��%m$jn�kA0Z�vjE?1�+քD|^��y]/����"l�\��R�.k۪ASO��Y�\ݢ߶���+�i��D�Q��Ng3�=<�Ls,�ڶ}BQ8��aa����؇��sF;���dr,v�?��;ޤ��(��wv�+��c��俟A�&�>���C�ʲ�k�M�D�[���Y3n|��=\���H4y1�&��k����ʢ���5��糶�'v21Z��d"9����}M�Q���򻒪��&.�������n�5��KyA�@�.��O���]�@����Qm<�!�-Ĥ�̧	����h�eCTb��Gc�T=���k3 �_n=%�J~���z�5�}$*r�؅A�=L�����K����IJ�ٖ����:�2+�x:�썹��c���o�.I�|z�W�R��p��"�<���4_hR:���W�,!��P�m���*����w\�=�6ٹ���"����P+bW��LJB[F�8[:����T7OK�]shv҆� ���[�mw<��g��4��6�f�Yn?I�4��e2(��(DE�QU���H%M�v��b�w.s��q�h���DN�u_@,��i�r�JNk�(�g��y��J:$z^��ZL��r�`r�T⿉�匂19*ۙ�c�ʗ����^n�V���i�j杰�n�ԫ��fݲɣ� ��!�Nkƙe1Ӿ4���W��u=(�x*Ų˲�I)A�h4����n����@Hk3�{i�=�p��������]�|ͤϵ�a�/�Bq�\�]5jja&�o5�l�=���gn#�Z�&�Dj ��gmRD�����Nę�����#���j �+(ИY��ʮ@@:u6I�9�RDn:���Q����w���1�X0�"V��ļ���̈O�����=��!�4a��<Fbi��z$�a�7	�-/c�*��	+g��q#���/� +sV1����ssyc�l ;���S�C! A������Ig/���R ��1&?#h{��.�.- �<����{\r��+��%���i���c[�F�	<�`���'��KN��Bpww��w��y����f�ݧϩS��j�sc��h�CP���2g�����7"]�8]%o���Sj_6�&H�%�P�_`y�k�=�@='O����Z*Z�� Ś�g2P�{�5v.$~a���2�^�m�f�������g��Y����F �U�K3_���������$|]�-�Tj���
WM�kd�|����";�o/�H�~9������f���o���L�6L�H;yj_��\�-q�k�j<����`����m�`�<���3������;���rY�M�Pn�6a[9XFE�ޙo�]�u�o)�] �Aq���{�+�� v(�ܜ���%���}��!oc���������WZ'�z|���zC֖�Ҝ�"�zϛ����·:��A�tjmev��Ӫ�����_`�)����� ���F�^_->��Es�G���~���$��˖�)2!�F��;�dZ��9�̭QY0���<����T�<���׵��D�ї�;��rх�HGv( �I���a	�YY�2��+�K��x�驋�����I�JӜ�^"[�?��w޿�cN�Y�upH4� �/(q�V�����`�hqPd�캫�=ws�~2�>-�}�����rQ��S�LL���Q��*ۇ�U�vd���㶋�p�U0sJ�*�,�����F��f(�a�]5�6��7�J���#��W�w�H=:m#��ߊ�h-�-J�JW��,��H�-�̲4o�F)	J�j(Ye��zj�����!��s،E���f�H]�T�o",�Tf5�ƞ8C���D|����s��Iy�w��q�:#� ,��o�Pw�^���ퟗ�����j>�t�t�v�[y�E��8N_��ܿ*� �% n]����ڬ:��eD�m&�UG۫�LB�{�:؎����$���Q�zw%&T�m����K�~�
�x�q6���ׯ����+��� u�xLĹJ�*O��4{lU]Nd�aF��!\�7"�T��6M{o��à�m;��c�1%~ke��x-
�b��K����������F3V"x~�i�x�:�	���mp�$6б����P�	ެ�z��C�X�cZ}���*�d���n�.g~�K0����,�I^�8����=���3h
zt�.�jn��n��֦3�jtMAf��u�e��b�H9�V��7Ȅ�*e��'������̑�=��l�n�*>�L�>�L�d�<V����~ɥ�Xl�w�� �(�Π=���FY���ӥ|yo�b��里k3Y
�زq�_��7{~��8�f�\�;�ǻ�]��C���|L�YK��贉k<ɪ��I�, ���~�M��s~�~�4��ϋ�TetY���Y���6:C�ݶ�����?�?kx�0��h/�*n8��Kw1�E��m���g��˪A��g�/|���m��C���H0��!t)�qp�VEm��Kd�v�a�싟�	��&��
��J:�zz���5SH�ns���>����V_�C<7�����;�Ef掠�H��u�)�ej���,6��v	��k_^����r b{�u��/��9�%쿛��M��5Vm�h��"i��x��(�:C�i��.ج]+��%?|��V\�]@��~�a�f�3�w�Z��ۃS��'�BǙ��gi�l�������j�"�Q[�Ȝ4��\/f3�����q�-�	Y @4>��&�0�{�>_���{����h,���y��m7��������7vh��U�R��J�����ui� ����Ͼ���9}$7v�@3�J��oZ3WϢNe��خm��}8e�ei��g/��FDq���彔���/M}D�@L �}&��������_��BQ����SJ06�FU�ǌ�2��J����'j���o>�e�7�Һ��6��Ԅ'��ɯ�Z�疋*}6��g+С��x~�u���.�j	��/��i�s�opH�o����?OưEkJW/����I\�u�S��[��t/�U�<DW��tls���^����߿.��)e�2�I{q���{#H�:�1R
r�GA�%��Z5E��}z[���lj������]���JN����ifϣCH��͓ݾ`�d�w�kt�6��<�#��e�HAUCd^��I�*	�,�'�E�]�/+�7�ή�ë2U0ɕ*�����&$"���e�%���f\ݦ����Url&��'?xM�/4^m�\9� uA��p���#����Ύ��'���2����W�˃��>�D`�ZF1.g5��ӽSz�Oq53�l�%�c��C�:,���@PevL����(��PDjPI�e�cH{� ��9��L��l�d8��������r�MUm1��Q.�z���q�?La���+������m����dPk��Ul������d��k%�ZJ{��������Z��6����D��O\�1F�[�G�}���y�ƽk��8��%��Ɍ�#<t�N�����k�z��_F��^Ʌ�*�o�A�w�-	=޿��&z��R\��"Ɵ�v�\RQ�ϛhQ�GS'`�QmG��T��������������)�#I�`�=$���I�;����x ��d��!���,�ӛm}u!k�T|�|�;z����f0f�޽Ǟ�s���&2�UZ�G�R��8����-��
'7�}>3uVG��Ċ��z7Z���
�Φ_��$D�Zr��4H"a3�g؊�8��z�G|di8�+f�L�AH��<�ag����]k��Q�OX�aG:j�p�:D���iQi?������e_�a���VB�a�ΐ]��;<9��7H��9~Qn��y��G����,�`�文�����r��:)��ר�a;��۴��9��jq�L����n��v6j���g����O��L��i����|�i�{³��膲�}�j�F`ϛ~�q�M����<����܀�l;��E��!��yCz����JD�|���G(C6Kc%���gΟ��׺��܋�����N���+�O늞7ɪ��[$!����%��>5���q�;�9E�G�o-&���m�"��"K��_o���x��d~��������� .d�l��Iծv��X��R���������2a�X���1�"��T��d�	!yr�j�ɷsN�rj�e�]�LH����v��h��Z�_7�7Tt�g��I�4:82�k���(T)[T�)˴nv�����������<U�?C�g�K�[�~@7
l'���N�6��t�NciG�F�g����R�B�f-�%-�\��+�d�m�.��$��@�5�Ě[)�X��v>����h]��=���- fB�5}�;	�<ͶcDO�+Wv-��:.e�R��`M3�l�j�OxF*#������V���\EiZW��屄_-˻�T�H��]2�ա�_�����_{��@���
�J������X�e�x���D3{AU��daI}?Wň�������*�f溒�G��}J�����|n�Ͳ�<G��)���U�Ōʖi`TEq�3������������pg� w⟿c��G��&Ï�/�A�*3�j����j�[;)��1��
>�4����ǨO�Z!�a������t��-RS�7�l
K"��@�?�I�.B�}�d<�������������&�r�a#ʊ�B�ޘf�y�c�W�BZ��aweu�-�#�4�Ś�4�~>�8��H�dg���q��O������U��>��ʶ��W�����63�^��t�C��v�~���u�b�uG��e+=<��<����V�n���dlZ���y�%7|��8�`�V#�M���"����߬�$�[�P�mz�Qy�8��_��BM��ww��������,����vS7�R�=�XcG&N�E��4=YqT6 �ɺ�p�ヱf�Q2��r���\���T,<H1��U�pd�+��%��XtAV[�C|�e�۴&eND�~�śC{��"'|����r�B��oF-�G˗n�(&�e��S�Gט��Ù������S��Ef9�E>�}9���vv�P�O4�<��Bo����C�n��K+x��qp9JEt�-�cy��	�C�U<����L�E���Z�s�E���j�I���Y�U4�ˍ����S�EZQ��C7ꌂ� y�D6 �4��,k�D$^o]@�+��IB���,��o�^Xz���[}u�a+��@�g�Km`_����ɝƭ�wJ�+�	E=�)���$��뢊s���p�q���H�* ���}�7�{v��.��i�Aכu�8�L����������ߊL;�6|B����bSW4�w�P?�֚����魖]�zg�x�m��3ӘQf[T�5�AI߷���h�w��9��b4d�n����{��\��z`K��7�cz�ak�^-̪h�\��*z�򏣻劮r�sF#}��}�Ie[�����Y�<�zR�b�������S��x���?��n���܂�l�:�~9z�J.��j��o���JL�V���*|�}%�����xفv�r7^w�����(Ö�=�\�Y��W̧��[ĭ�Դ*p�֋�>�W4X�a��g$�lMJ=�o7�Z��SM߭i9[�r�"Ӟ�]1?�<!�GZ��}O�Cb�S�40x5�ɚbFY%��'���&��Q}�rۃ�R��D���槿et�~(<&��ڥ��6�6�~{��z[��I�m'��c.,����bW��S��(*6n�Q���������dmw.?��[�c!"!�uS��T�K�YZ_�ݘ�O�pF����y�o{	:2�_�"R��i>�\gm:l���8�b}qz15bv~u>�M��|���|��aJ{����1h���vB�9��� �nhয[=���k�p$Dv�2���{��N�-P�2x��f��`���_i��U����גv�l�VM�g=c�h�őP�1�����_y}$��$�%1¶�O�������|o�u��:����lv9W� AuH��h.A�_1]X׻��O4d���*�N/��p�)C���SN�~�����CAt�#�sM��N��p�a����l���>����i�-��S�:��x�|�lu���D��w����~�|-�b��u4�g��0X���n�a�Qr-����C���(�����Hh.N����=�i�>b.�	A�}ĞU�uw�+<[�^���홗�G5'���7O$���W|����I�WS�����J�҄l%�}2ha�4���/W��Ƿ.�.Վ��:�y��`��]~g�Hjb��ԾMRX�o�2�l��ʐ�a���\%k2uy����|��� ���F_���45սO9~���#�eȱ����bj�D�8~h��0��7�a+��xnC�I�������Unu�Չ��m�ʻ���K3�:ݍ q|�/�z�����ˡCv����TZ��ՏӱP�4FZ�;o�WV���҅FQ?��V3��巈�XP�N�y�^//��^u�fus:����F]Z��~"TH�笐A�o�]:p�c[+�S�0	�����p�����;P@�J�G)���.���_��Z�^b��޾�t��a'��m-��]��M@����W�!� �̟�rNcl���L�}'�NrT����9WP{_�����&����������8�Vw�����&�Y��DTE�!$4�[���|l)8�O��<�R�mΓ����(��Xm������S�E�o���ݟ�Z�Wm��~�d�)�[�6��G�%4y���x�6AQn�;��������!`��i�S|���A��gpGVhV�vG�ͭ:s����Aק��;s[���?%�+%ۡV����g��_P�sJy�s$~��M��{T�L����qy��D`P���I'^%��x��Ϗ��<h�Ə��R�]�-*[1a��E:��Q��H��i���j�SJMW/�M�DE �2}�R%���)��֨��4<�(b��4�������)��Xgց��}ZQ��C���~��5?)n���zC����Tg;����9P�Y��׺��ų���ctj-�q�d�}C֖;�n����ݗ���^ͭ5-���8���3I�p��_ۀi�p���#�lw���$�w&��n���~&$O��M��ޛ�j�'�&��dD�{�u��}0�&� �������4HI��T,���&�`�GF<�9��:aK�R���M�B��t;d���c��z�񏥙�v�����;�TΖeN8��e_�Q��}��"�Hn���S#^k˔3��T�ku�dF���:1�/ͥ��&b��כq!j��`z#��k�~,� ��74�R6DDL�%��[�|8��Q��M"zT�k�?S���K"�7ܷoJ��[��3f5F�RJN4�s�7�a�5�)pE����\Pr����O�5��b+��ۏ	��K�9�O�]�Jj6��k*LB�F������'Vʽ�,�5A�{y�j���"�E���h�9S����	�U��9�M@����sU�@ߣ�`*�|�u��!����Ϙ�E"�h���Hw�� �
U�+}� ��L�@���"p�ٔGe�@�^��"�/!�/�on�=բ�������<�,栦��,�Ios�!��x�fFqV!(��q�u�Ջ���Ε(��[I�0�����1����ԗRR)�kS��cu�
��Ȕ�Y=J $O�Z-?_�H3V���]P`N7�1�V�Nu<|��;\�K��v�=C�����y�~>VXs�jʬΡ���}[%����� ���.?hS��ڊ��ۥ�7��3#���	d/ɮn=6z]Ŀ�	�M�A94e%� Α|�ݲ$L��唆��.K���*�V�WoG��:A�ǅȃ�]"�.�ס���R�(3V�z�q��F�;����ؿ�bG�����j�P�\��ڰE�4:�rn@).�L�N�L
���(��'P�)��y*�_Kp7B�g	����L	D9#�7��ƗE�~/��r��p��������>Je��Z�̦\	(ؽ�AR��&x.g,��&�*�ZvM/�������{>�G�H+�����I�� ��I�?kŃ�S�T�����AT����c*����n��}��s/ʜaG�Cn���#\D�(�3���뺘���&� ;�����tt���C��F4��Nەqur�.��ucP~B�wpk$��T��_˒@��"�nP�(�n�:*�3���p\���&H���%�d4����!8��4����N���m�����$TK�~�T�9l`eu���;�f7
}!��.(�X^��i&����~�{�k�QN'�l�3������+J9M����zz�Y.	j��z��On�B�$�Q�� ��B�a�:(���e]p����&��ܷM�ñ�?���H6�t�MFP��Ih��ʪ��Nr�=���|x6)��iȏ��~n�C A5���\�7V0��顦��.8xh~z͑VU�(E�_h7&5�G�P.%NyD�H��6$M"3�t��^p)�2�h];�X3lt����;�R�!���<���3&H� uPOǢ��s=Z���$��拿�Rh���!=�}� 3�(��l0җ
��W��hޟ����U�e,���+�K_kE����q��{����1��+{!.Li��y8t5o=:��Z��y�mo�چ�:"ZgX�?�s�������3�� ���?�Ǳ<K��o��^͊�����%�z�[���گt����/������;�b/���`j��ƒܼ��
ԣ F�������W�G�����8��]
�L{�4�
j�,#K�D	�����9O/*�kjs��/��*�ԁ�c�.rA�&�d�>xc4�����������>��?g♊����A)s�d�{�_$��\^Re`��qE���;�Sl��FD���𫍦��)8�k���ߢ�e��Z0cpnzF��*p�cӐ�Q��x����L�,��_�48���}�2m�7�=�\�7�&$%k�����@��Qm���#���\��q?���ka@�4B�AB"܊�h"�Z�J]E����,��:9M��_2i�x��lbL���h��Gt;�]�|:���Qw��[M9"�4狿��*���җ(D�![�����A ��$���J�LU>ex�׹���t��VK	�(���.5;|h�Q.���L劙�$H-9H�s�<T��帀R��ʬ�}��Dz�n+:�a5xpa��5�L$�� �C��
�W�ϒ(Dg�9�����DG�>�C�ty��_��z��ғnk���Q�rY�@�P��������h @�~� ����Q�g�.�9Qm��v�� ��]�z0I�`��XC'/�7�J��n��L�`S-�)��a3�	����F+}}�YemY� Ue���sR16����|���-^��V�`�|�O�v.��G�sX�<�`�مh}D'���Th x66	�v3��`H�)���8���K
����!�h��	ZNHYsC/��m��/�Xﰸ7���b6ɝm�4��x��\J��-<S���v*��������X��~-��.��%��D�Y��<X�$O���"�mT�b��#꽟Ӂ*�;�p�@u�K���B��[���]ˢ�.���[r�����o,�J�`ْ0Y�:gg#Z�_�3t�{9`I���^��������?Y<9�x>����1���
�92��H׷84��}�?.�J�(�������xp�q��76i_�H�ʽ������S3h��[L� �j�WG����õ�=U�u���h�{G��Ԋ�u	ae�/���;d��X����9|���Y�� ��U��q�/�2F�(��Xm��N7��-�Wy�{����tr��g�kb,�֚Ƶiz� Q����`@�{\�U���wx�גM%���v>I�d�/=����Ջ�oy	�o�5��٢����*�QT�G3Zw���'����7�2U}�qu�����smD6��cK���G�$�J0�VQ-����Ƴ1���6�\_���M��b.#�[�����'��$$,������>Ė A���ɇ&^RJ>�L�����Ȭ���g�+d��� ���ʌ.5�CX/-�1��N���5K�i9�4"b��V�ֵ���!�QL�����%�^����(���>�=^f��x2]�#���I���
��=��Jqf&�j�4K���m�U'� P�ؗե"$͓���?Ʉ -0<�-KY�M$��56H����������p �?���Wb��ݻ��+�м^;N�j|��H��x���X&�	:��"}�%_E�>��n�?j��8��&��H)[ �i�M���~e���E�4�Qd&��
<�Pw�Q��عV����(�C�$���XT����Js�e�ד��j�vx��B�[�LZh�^�T�����dyv Jx���OW��'��*��^6�K26l����|�{Odn��6�zs�Q tT��x8�J��nӐp��&:���9��n�&?.�:��p���� d<��J8TPR���.)�r�zFyO���@����[Q��*�'�T!Lڞn���ཿ�egQ��J�^Rz�;�~ĕ"q�_�o���Y�`5L>���`�S��^	���t�?27�LqGJ��������2j��DJ�G� !�I����˓�I��f��wn��倾>Ijo���M�
0ğ�Ʈ,��Z�4�XٳhmJ�V��7��Z�>A���	J"j�%���:S�,�@���'�۰�> �H]�e���n�Zf�"���৊
L˔�d��/��k���Z?Eo&2��L>wr>h� �8~36�dt���P1tXF(��I�3�C�K�ۥ�{�O���>q=z���Ķ_�M����ޢ������9��徊RިP�.B�^�ȩ�l-Yȼ��@��(Ǿv�LYy�F.�1d܈�⧀F���M�H�m.���ӈ�yu*�be a�	���H��iȀ�a�s�@��?�6ӳ�MP!w�8率�gc@%�2�g���*����8��i:]�r^��]�%FlB��ms��֘?�nu�y����V�'��� ���wz^p*;Pa��X�h(;!�Sh7[Yc����Y�H���P~	�ΎK|��L�_[Y?&ᯰ�"⩋RPZ�}��<[T��J(|�(څ	
�K~��!%��%В�=`27�IB|��)o� �:"@Ȃw����������j�V�õ�����膶@�*�/Ĭ�b�<�AU&���o�](W�T@!q�$ܯ�2An�S����7��ʴ*��T�Zf�����}�J��wu��Į2��M,��t��HJ:ǃ�]�yj�?��E��~FK��=6X�	�YD]����1c&�n�oS���Z����Sޯ���XԵ̆Y��2�C��Wq�߂}kI�U(d�a7�q��I��>oj�����Ta��z݀�-�D^��&Q�<��<�.�A�q�*_��	�S��$���h'�GP�$�4��������c��}�A6=F�[cL/,��_S��=K@n�+.���W�px�qt?�W_Z2����_�Pv-Jz'c$��0U&�!�'�\Y����a� (��Ν�A��1*���v��l/윎Z��?�A
���e.C�z�x�Ԅ��c����;Qs@u�77$�RR�t��U
�
>թUY�W�����_��O�nP��]�xT__r�~P��&� ��ݡ�o';�����( ��k�DiB(�I��0�#�K���q]�IF����������f'�#@⺷�j��ɤ�/�F/aD��q�v+cZ0�{��m��O�Hz�JVy)ԃ���D���(�����YkJ�,1(�!\�Y��ϓw�8��ä?:\J��"UQ.B����c|E��/��qj�X7t+��%��W�9�U�������iZ����{0!��ͧ�c�� ���M�P��ZA?�)Hfm^���ya7�"�(���W7K�}���♐��%�
��~�<j����2+u��Jө�kq���/d�/h�D��7\D��0�6�
���Tn|x��#�ݬ�0���T��#�	#��)P��ѺC�;��TE`��,@���X��v��xcu��Z4��;���=�]���iv�	�k
f^��{r�>�J�ܦ�w����4qX�o�q�y$�adF��d2F8Z����k��֝��l.GحLm�����$��G|��������l�e�`�Q��Hi<d��5A�U253�]QAB�z���A��2>	q �3nq���ϣ^��C�6@�ޓ$!�J�f�{��/}p�uֲpN!���C(��B)8Z�j�!�"|�P��-�7#$����#y%�zwZ-n<@�j���<7�>͛v��k�������a�}�q���췬�eA&�*R�BȀ���hx#tWI�DmS/�̄��M�R�`O��zx�U&���I�ފ�'H�bu�'"�|��YA@6M���Uix��2�� � xv�/hN8�o@���di��
��k�Φ����PW�,�^Tn��B�|(�}��3օfm{|�T���~���!ܸ\����W)�(X�{<4\�f7�+�d7VA�`&0#�����7B���J�LbO��;�{H}- ,ۏ@�d����2��v{�	s��d�[���j ��2����R�C���D��$!�~p
ղ<������j�x�� �fl4��4Y�E�b�A�*��%P�/ޞ��,��(�����B}:�[�F��/��HOp!�G/���t�n_����!,�����E�/��8���[y��VdN|����P�p(��ԋ�CQ��}����dD�3�?&�e,L�2�:�9�?�9Nؗ]o�|}���c�(�1��o���(r���^�R�a>�=^�B\���$����@�����r�\��<�畉� W/�y�Ro��0O��0�Se+BR�o�P�G	+UL��8�H�K�;�'��'k�=^뵫[Մ��(U�&�F���@��{:��d$�8�qI4%-�ԌhwP��f2�b�956�?�h:��!�2�@W�Mu@?#��L�b��_V�И��Z�ia��q�ڇפ�Q6+���[}��	#4E��B�(�j�m���<c��mOߵJ��=���9m�C
e���7��h�q"�$w���X�P�e?W�(���kY�O.D���~BVܵ���O�L7tq��s=�'�xCTz�/����
�?�WR5���A
s���������OU^����I��R��_�_���f݇1s���Z	{[رbK�D�����Ǳ���()��40������+�፲���N?��v#Y��FSVA�`+���|?k�9[�%��:��H��h�c��и���;X���*��9�?V �^�]";�n���0�bx��'��}e�[���:�UI�-��$���}\��t�� ;�k?/x�{!f;�C|��)�¤Djj�݁���#W���/�`Π�Pb^5>������!�]br���VfC�"�c�O���fG͹i���7kY1�r ����A���(�h�K�qҧ��N%��ۗ%Q�x�)к|�ڛ�*Hg���N��3��m����PK��"R(�n&���48��\}�2�W�Z�jW�� ��������&@s������\p�����'D͉r��2�)�<�-�f��]����x�ĕ��pȸ���i5]Hr���e�M��%��EoTkL�������PPhv��Xy!�Vc�ة���'�-�a�"y�zp�R�M�f���̬I���[i�+ߩ�Yf,�71����K�5�>`�����|����P�*�����_rXȡ &"oAL󳖂60⤭�֬J�@:����ޅ:�w���`�|:�[�~e�E�P�_�s�����c�0���;�3˽��N���[�����xY/ ��C���.��;D2�ܗ����8)�-��+��B������V	-��C�V�G>��2���6����Q���2Q~ۇ��Z��z��Io_��pl��.�b�VC,J�%���Iqf��+�򒙓��1k�ζro��0�l�bD��ޟ�g��&��+	ƹy�oG�������]s��PMT,��p\��to6K ~�?�����Z�u�N�H�O��&�l%����:�3>�������ʬ��������I��*����R���tI�^����Q_��~�$K�$>����|���������"?���6M�ĭ�GD���Vtm
��V�6#�B�No�N���;I�@{"��J�%O/�j�cnF;T.�q�e�E0��i�@u�k@�{�
��o,2���θF�f��s4eD�'�&��"`J>6�Bb	QOn�,>�NR7h@k�h�A�d��������QVAbe�i\��c �*� g����:H�L��ۙ�d;'�6S�C��px���E���|��V�$�GE$���A�2va4 ��1-����@� ���(�Ҫ�7z�䠁!�(@����>jK�c����H��ȝ�~L�:,f��s��>��� fV5ܭ����X��@���¾#~�qH�g�z����X�pй�r�������� xIN��).���ݡWst]� '��LZ�p��e� |���%^G�>]P��!���t�;��q2�|��(�ɍa���0S;."�y�k��*�c�婁[��c��t��H~���������M���{T&M�K�)��y�&���Sd��|$���{�1���c��/-�S�t��/N����laU�//�����O�;� z�)8{(�n$ͦ$��5�P+�#Z�k�����׉�ѻ�gm��j��ʷYs<��x��ϳ\�Ý����q=��jF�l�߈��_cSl�Ai��c�Hm�t�U��~��:��M4|����o����ř�r��H�f�_�NY�HZ��^�H�Į����ĭ�f���&@>�5�z:hR6G&�%
��
���LY�[� ��V$g�U����&!b��[�X
z.#,LVu�VQt��u؉k (���[oiw�}[������鲞����@z@��'w*.*�ԟ!�x*�hdoct����p�(-��nb�*�)�ko�O�v�o� �#�3�cv������j�'`v�cz�N�=״A��+�ol�C�'�N¦��9��d�����p
N(�&�����ɔ�@}�l�t��j��n/MZ�����-�D�=��A�;^�8�W�^�U�S6k�j�p�V3�>#�ldC1gc�.�p
N�-d��
@�a�v�z������c����fQt��N����E-�i�K�;�>��(J}�R����2UL*D,�C�o���o��K8l�-e06/�A���8q(�]�4G�!��VN����t�
����H g��}��8j���P�tg����(�i�p8�	�{k��2D%��2��%��q||�s��Ǫ��iXK-k!NƆ̒Y����q�"xUP��M�Q,�^�kϛ1u� �д)�,�r��	6�FQ����$q*� ��_� 1���)�?��uD�X�?;˔�(�p���XG�Ƿ�=���L�,���APP��g���_!t�=h7��9oP-��z��3����޾���C{E0=���̆-���?C�6�N��V�,�8g�.#�o�>8��SGCo��k2:Qo�ͳ��/.����[zX�G��A	���x.�K����΄���Q�X+���{#��@&p���τXVAko���]b亍��d�%8���,�������U"r��1CI����(B��%�<~i�؀"���>�Xd $�R�Z3t\l��&�s�־�_�K�Z��rg�[�#T�ex����a4�a���9	�2�$��ʠo������}�4<-��"�x����G���mi|g+�3F{���C����B�*Kp%`����>q��2�P��Z݅�ޚ��0Pր���zD�_X�_�S!�ޮ�.F1 "��ᢶ���#�nɿ�.}�H��R�=�P8f�) ��,���}����u����?��V�̎���Nm�n�9��[	�� 珆�Nu��.>��Ax�ϵ�g�����:<��I�Ezj�Q�{�N=���o����A�o?�x���i�-�Ȼ��]&˶7QE��e����s�����=b�I��Ό]%�j5��l�zL�����p�.cv�̫R��jُ��,��"hT����a(���R�C��1WZ�~�Q��	őFt<����|ԇ�(��X4�g� w��	+-Gq1r1c�Y	�,�*��>�a�̰P��(�ۻ���=�PtR���1�i���&�g�G��$�PJ6�Sg|�:���,�|�CC>���iM	)Z���Ƈ�W��h����j���Jc�xk��}�8�׼�T�G)F���P���b�X>�g���)����5۝pa�������(��Y�'$
!T��"���B�mΟޯ|�i�Ò��~��L��8���PX�z�\��Ì;�=O�4�;͓��:����#�#��Fe���M��r+�o��ʹ�*0׫���"�#}@zm���k@����:&�֟-xGC>��y݌}�6��5�w�c�^|��S'�kA��<�9�1C+�.���'�W-���,���Ycq�[���V�S����j���G72m܆�NqÜ}�8*i��g��t���#�o6�$��ߥ�ҿ�v|'����J)%��ul\nٛ���ei��I��Ό���n��G˗:�Ai�#�f������}*��!-��w����ާv_i��q���v����GG5�5�>mΞ��K�?7��{#N"����<��E^.���;&��<�-ԌVvl�PM��&��S�����˨~��d0������֕`4*3�2F��ʤ�mv�aN��
�#9��7����*��X�F�M¯@C�&�iA'��j̝�s��^�|�{�CvC�=|s��+|�]�;_>_O&J�Z>�5�&�F���nH�2��p}<�|1��{��&����|I��3H�!��y�|�cM�l��JlYl�D�3ϔ��ji������;;h(��W+1��� PK   �C]Yz�� 5& ( /   images/aa32f2d7-3103-4396-8365-58a51d23b1a5.png|�x&M�6M0�m۶m'۶�L���L&�۶�ض}������g����]իj�����V]W��QJ
���q�����KK�����B��mАG��W��^@]T$E@���N�v�̴����Ah��� ��( ��@� �8 ��e��h�����>(տ1`�Z���<�
��_��(R����d�ifkg���L���@������w"�_hk}>����O=P�|���n�G�������������������ęͬ��QJ���

���^o���%/�c�`�`d�`l��i���{����kڙ�y��ڻ�x������g����_W~-y%"Qg3"&&��DDD|Φ�<*b�����X��:�02zxx0x�288[02sss32�0����Eлxٻy�ۻ����ꈙ��8[9�Z9���72vps�'!�7�?�2���H�.����	2��adf`b��hg�<���$W+��C�<�A�/�?w�����3�w�;66>����2�������ߙZ�+���xD���I05[��-���'�0�[��1zfz&n���1z&.&��&����!�7iL�\��*�<O6�������7�+��������?� �����02���1������_.u{+W�S����di��j�_*:[��M�������c����#��c1�{	|��X�s?
|?�E�V�=-^v���^f������M"��J���~f�������l�s^�MZ�/���lz�^nT��IB	R�#�HI�6�L�uп|zu�{{˫�1h�f�le�o|<<m8^�>����G�����(�/���nL�T�z��6���T��>�|^�x�t�\>�&Ci���b�kpo�Y�J�Z��z���k/'v/]�9�9$����,٪W��j�-���V.Z���F.��a�\`�^T��pd-���u�rv�ZQ`�)�%D1�n�u	�,Y�6��Μ���� ��	��)]ReK�~��Q�U��H�-���VhX�N#���ѿ*WkT-Z���-�ٿv�b��]\,~��R������?����l؟�~�=E��:��>��?��a��yBC�"�|r]k��T�ky��T�pk��-ث=�S��;����J=�蓶�ݡ�7��E�4�{��	+S>����?˷��"�`.`������}���M�R���9D��X����?�nT�?a~+��\�@�bPO�F�?�.oG]�|z7[��AH�w�[/S\N�X<[�N�P�Z��e�nƁ����i7Cbl�������m�]r�L�
eJd���z�"۠[p��p����D�V��������x-x�zj4"�,�r/'�0�&/��r?��p;=�T�%� l����L�lR�p)��m�4� �C�ˮ��u!q��sZ9��?A�'�(��o�ƪOb@����A��������ζ�-v�Ś7ut�#q<��rA���B�Œ�Ώk�.�o�4?+>��ˍH��:����!�p���A]f��ɱ`�b��;҃6���BC��!M`�#<:^|<�}1Y�J�\D�'r�Jm���fv�<�˖woK�u
9 i{���>�'�]�������|�mu��s�:��u�`Q�U�j"(�b�hH�Ի@����Ϧ�����Bٞ-���Hr⑴G�����F7������K��{�a�:Kv ��S�� ��-(y�n2=�T1�B���MJUMK0)=�p���kE��2�^Aj�l����̖Z�H
W�����p���0���1��`ؿ6[	��xu#�޹��~c�OI �rQ��Vt�?V�$��ܠĪ�gE�	:��v3����x��TZ�!���~��n�f3�	�m���)쐲�r6}Q����uL0ϗp`�;ms��s��k��y�~�Z�؅�v���6A��H�xyK�Қ�H��*`�5�W�!�u�n^Q���$����ǎ���ǕՂ A��I̢��܆H�qu�dʌ4�8q��<?Mr�1��$>`<�?1�*WKz#5��8�����[!��X���#�6u��$(��c�y�ǵ�9�f�=�#aB�y�@_�.I��
�̷'`��'D|.*�a����֞��p�+p�k4o��[J���2=�$��a�h��ͥ
-���a{���)V��!��pB�L��.�2�!DMޫ\+���G��8-��\�����T��_~;Q�3�rA`�1��#���t�pz�i�����u(�8j[�(x��+���zSx���ݧZ��F�e��cma�B�?���G��7Df�����k�WL5q��X��-+ݘ�_�І�탋��F�6(8���C&��cD����D|Dߙ^�ªȮ6z�l}Н�$Z�y^"J���֝��d#���'�r�evM8p�}
R*ol���K.�����L��2�Z�zIKE�5p�m
I�S�U�܋k��n�����$��+5�kP��_~���E_8�k<AKH�b'`P/Z�HJ�4Cd���bX�a q:P�;P��a8��
�S_H�{�~װ�;�y�
�_��3��,sN��NB�zCbGJ�����*BpkcS�ŵ8%�S�ohL����U+b�=G5��#Q�-y)��=c�q��"����BR���Q�b
G0�X;�m^}�#�8fwq��\�M����>$�Q�%��#^f>S�Ī�z�a*r�1^��4e���&EK9p�]����d:hc����Kn�`Y�̸TŠ;`3��x�	�IX.�6&!$B��8�ge)))SC�?!��i�F��:TQʩĲ��\_�L���xДb��cۋ���� M��[6U����2�D����b�s���g,S�����EB��}Fh`{ Ro�Ӄ�@k�/]�U�t!��hG^�h(�g��R ���� ��c��~9��oNt	����u\��r��)�r{5:v�E�w.E��_�*Ԇ)KF�%dJ�#c��J嬠�S?�0J�jA7_�k�,�@���i��y0�*pkU�mc�3r���֣A�
�����B;�DT�
������ȱ��ٵ-epls��H(O%��΅��2#�+5Oq�*�
��hY��s���A� dfyө�����G%�	EJ� 	7ʛ�FN�I�Lp���uI��p�yޖ��o.;f$c4�RF!2S�\��.��h�4���j�(�1��M�7E���%�Yl0�qN����J����X���lO�N�e�V�C����^�ɰq���h�c8�1�)N�-T)�V�6�Ta7���M���� Kg��VbN�K�н&��ą(����� *r@XMi}���a����$���i���o��X�����^�2�z�p���湑	�PE`c�Z6y���I���y��G�g��.�d\cF���!W�g�d� ��8�D�[��w��{��&�<��(�s����HDޅ����\��y9e-�G�О��ɉ2�HEF 'Q҅�\��]���!��҂�(��-�C��Ȧ�\FW(Z��ds��I]�^����gFƀS7'������gWl��nfp#t�2ڹ0\�e 1Y�`'�x78�]N��e�-U�IuȽ�`�RyM�D�Y�嗈�Hߩ�|�6���j����*e1} �;��Yvm���+�w��C9ܠwҢ�v(��E�-Y��^��� o z��7�M��"��<��B� *q�ԭ����Úaw"�͕YQ���TR&�ŞE�U  �[>eR��=���F�/PkHt]�I��hoE�/�-o�'n��oe������&b�X�Ʒ�?���m�vA��*�ٰ��!�8���i���!�Q�,g����l���E�\2�1N؆�fˠ��`Bd�֊c��6y�Ɓlq.r��(�6�wv~�
q,��Fu��❠��	o�� ���m��3~�r�9�^�'�9�G�*-\��[�f��dr�Z���
1����O�����֨o��\�Ğ�#U��c]�-����TB��슡@X�R����5"߄���M[�.�Ԁ|��}�]�v��C��,a�$�t>6Z$!�]*3�>=��t1��I6@��x@�"��v���0/�7~U�fB��~�¨ �f����I�]����~ʎk�b�Цb���&ɢ)�2&Է��Ԯb���d��^��K��/��x�
�pۚz�h��վn����Y�;�L�[#K�l��O����cN��y�]��UCC��F$�G�i�2�Q��v��X����w��6�*2�
�o��W�
 ��e�ۏSn�5�,)8�ț5���df�W��q��F���EN:������m!�|���|�>���';�k?�=�X�E">)����K�f䡐�`�E!,h}��(7��,��|���iX�g�	����0vo[�׀���޼Iq	!��Uc� �EI�Y|)%4�<c6�|�LI����)���b~|�R��l+��c��<H6�h�[�x�A�7.�
e9
D�u���k�.-�8f&�q��
}x�tg��W�U��qj`�fa޷��a[�f�̩A?����1�ic�\����^1o���^?�1?m�\�u��S=dk%���(g-M�@��,�C�O����X����^d��EVi�rh�բ޹�*ȼ6���Ȝъ`]�A�i	����v8'I��>��c�����"���rh�/ڛ�C�5�1H���B�OVU�:�����$pX#�8U�E�j{��[�����ez�n�!jT����p͞r�:u�fm�aI.D���ٍ�X��Ke��qn
W崃�B_f��qq�F�lɛ�t��bb�lٱP\V��¶��Ƞ�ͱ�%݈�zv"l��������k3��z������>X"�?u������[�~4�o˅�w�	/�J�.�h���0��%��>�e��D�A�ؘ3�t�P��y�:�T1;{�����UfE��{��Qv�g젉���u�k��?��?�j�k<q�2�_�b�$��5e9��r͉0��!lY�@����^\�W���}���1Dhf0c?�~�2!����/�h���`����h=X��ؓc@��͋���Z�㺘�b�H$?�	7Z~E��;����-t�l;�e��,���JI�{g��,}1�Z5{�yd�N��Bj$�I8fU�T�;BR����h��O���fe�V�<�kW�}�v�vH���b�Srf%�q�f��Q��OU���	�;|��DD����ʄ(����b�1��:���*U�<$R�āך{�Ukk.��g$���v}�y�ـ�Y���䚵�hƕ�]r�ƻpw
^{X��śQh���U���W�0*�\�c:n��/K�砿������Iv��\��'N�^h$P�/=n �0���v��K}�ye������+��k����O(��|L�rbs�������)^�z�}�1 9
I���	��KN2��~�W����	I�ʎ��+A�<��
y��j�o_���TѡM����~�5�����^YV����f�$L�t�]o�k(-f�@�|0!�W��yO�� ,�**�bG�_�Ա˺Tms��i5*�aF��i���q��?�f�4�s�ڌ�'un���;�|��֍�ϟzm��\�g�r��r�����'f��ɋ�e�n�Wk�u˽��s��<��rqu��H���_��l��R��� �isf$[�#�qQ��h����[���zQ"�f����=ȿ�Y���r��3��UR�n-O��2�+���z� sݤhyM�)=A�ګ�!8%�H��y\�y!,	?`/t�4�*��2�.M�AIZ�MBQBBu�Z#�E� y�G.�l?�Q�z!!�^:���7Y��JH5n��K��T̷֭�=1-��Ek��H��	[I�f�w$���f��T�ȗo�f�B�$R����u������ZF�׆3?\�Mu�1J{�	j�ªłF��#$b��@b�*z\�F7��V)T�_;lpL7yl|	D��U���zg�� �gmޝ�(~ƚLw�O�­�\�$�w��lJӯ=W��A�5����/�=�x�*W���+Kaqm� :�nHh'��v�vATk��1���>}^w`�x)�|�Z�8;����f�p�ڪp��u��ɪs�����}�Y���{�3�����*@eP8|��	�l��O���
S�
�W�-��g,;.�Jzv�Q��{���"b�UΜw�{/Ò�ƷA����%i��gʊ������H��ֈ�iSdg�Ts6�aE�4�\���QR�*SW����P�/�����Țʈ���.o�1���ʔ�ӊPGġ�p.���N�����)�ĥ��x��O��wU�h�X%;|!d�q�ݹЋO�b��l�c�XT��֛��}'7:<��x�uܽ��h�F�Rnuf�1��A�����
�e� �>Ӊf%U�ʮ��#��tz��fE�!ƌ��'&/���
ٟ M�z2J�:�ۧ@����oŸ�f����Y;�����:DY<jW!ֆj�` xO��M��qM��vW�f�-G���d�ͽ�(�[Wk:.�f���<p%�rB!���¢��A��sՙltD����q�F�N��F����/����W�����ӓ�R/d�l�
�����J�����
4-��;A�����|{�{���B^��="_�x͓E����q�G��������]��s�(8���N���b���'��s�&@,Mo'���fI�%'>!�d�da��읣�p ������_�}��׼������q�7�o�%�;s�yH��x*(��t��[$d`�p�z�=�_�!����^���MTө�	�:�0�o|��=U2.�?[�f��,�.��g�P�������6:j0/����"�؉�4����}�������Y��g�<TJX����h��J4=T�fU����O/��*�1y.�hZ���ͩ
eW��y ����+W��yb�����(���@�
��;�;��ee�}n�4�b�k�c?ѡu�.55��ʪ�X���71фu�3ؾ{�"�0,�,ת�)�^���HRO�|�ԁŔ{ȀIx���S3-&���9�&\$��d�y[�����3��o��*n�m����d�?�(1�"d&�@!r4_��Fz-S�_���>�Z�ߏ1�q~�>T��ڔة6�̑Y��.�,�{��Kd?��d��،���it���Ϳ����z;�vC�G���>(\��|��h�MX	����U0.NVT��J�	x��#�5"!R�`IM�H�"4 };��̥�D)�r����&�{tM;Ir�w�:1��������gJ���i��kh�������8|���7����p��z�F���m8>з[~��C;v�w$�ޔ XgA*ԍ_$d��eu�9�uN�)��Ѵ����"�?�)h�7��a������eF2������y����ZX@�A����j��+d����Ɓn��v���Rլ�ΰ��F��Lm6��H,0�V@1�n��H ��)ُ�i)��ԕ�
�⹅�������LA��j"长����IPP����GH�ib�x��y���~.���aߩ���귬��^_����+l��tOh.�m,�ɐ�>�N�m`ʶ��r���m��v��e� k�(��=��;�
f�X����>�)yG�APG�h��Z�=��&���ֹ��Zw��NA�t<_���n�;�#��n��ލ����_R�z��ʸky����#���~W���N6�L��O�a؃Y����k�].�i�ɕ�=�ױ��u�Vb[�d��,���B��æ�f���k����G������Ɯ�%�O�k�VF�.�,ß�l�ڭ�?����ME�/6�F��}.?&���=�o������[g�v�Y�<>�e�;9Rq/V�q�l�#l ����&d&��;מ{����Y����R����q�dʍ��y��?�?.��<"�á�ާ�Q^R.������6C��|_n]`]�S��J� ]�'��q���{���x;��Sͼ�#�oY�>��7�p𛲢>�4�r/�]��^mv~��J�ZG������{���=����4���m7o"��H�����x'��D�I���T�Ÿ��?q̉�*ӥ�.�{��+Ĳ~jK����X YXe�3�
1�1z�Wh�p��*";��Q�@�Y�U�9f�~���M����@�~�������T;���B�����F�"��'����{x%5)������raF6c�d`A�qF��8�E���n�����wW`>��(i������c_���!1�:F��Ȏ���D�r\F!�����ѐ�7Z�6�gq;�-���ؼ�������f~���U���t����- ����h˝j�bc�5�p[5~�{�K�ׇ$��\^ć������$7L ;�Q!����u��`�6��Q0|�P���$�|����ϺY�h'`\��[���d
�l��Bpw���,�
"]G�����鱺g0'�\@�o�����v�w�e[���99p^ZS��[)q�H��J|���)�	Ƌ���;��`���N���4�cz��8E<��H�$R�i�� �q�D[�J����!�2��	� ���C��b��`✦�K��M��t߅�Z�n3}�h�Qo�q��c4����"�0g����,X�]#����^ݒh}�J���ҫ:2��a
!���ZtˡZ��	���q��f@3���pl7��Ho�>4	�,�s�E�)��%�2�4Ă�����M	������oϥu+�(���·(/��Q�g��� ;�(/ƲD��(���vɅ&i�ZX�ihi�
�$�+G����bXn�kT8+{�|^P%���eX�K�P~���$N7���_�����Dc���K�?���gW]4��~,�k��D����Վϧ�k�c����]���{��d��|١����/���F(�P�9bO(����Q,���׈+��Z	(����)�Bl��ܘ|+
��x��M��+|�ݺ)<#�	@��p���H�D���%��'�:گ��w��)��-N��^0��A�/����A+��̔8�<;�Li|`�%	p�p81a�v63u=�y�lI�<��AB��t�k	� z�mL��瀆U�5�P����(��~�����y�3q%Qy�3��ʪ��KSR]�&��g:*2�^�b��F7!�QL-��V�uςw��[]X��-e�ih�_O��_\�Z�����"kS5�7=dBD��D�:^�"�UwX�1��%�������g�Q��L�w�Ƿ�ϔ��Eo��$�T,r�Ua4(�T�I�5�]��2���C݊m��Ty�������!z[\#|��J7���F�N�BV7��`rU_eTFK�
׷�]�^�$zS��a���z��������eΔ
	�VAFІ�v�$�C�T��Σ�	ur�ބ������U՝S~Sn��°r��������'�b�$��&) ��Z�M�V.����&����(a��+N~�b�$�Q�N�AP��ʀ�$��R'\�YҬ�M�#mI<�� yWTs��R�:n��Cw�B����I���ӹ\X+L���UU��)��((旀�}f�����9Y
���~��v��@�A���.նpF�V����,T1��k�푶��JA�����5|��fh��U9š�0tMt���o�".?K֋8a����x���^a\a��ǆu��+�H���H/�
KG=_^�����E�XVu���L��=�Ecg,�D�l�v����2L�#ό�>yqcRB��_wFl�1����B�b��Tʥ�M��q���~Z#��� �!�<�����b0s[�,g� ��5�e{}z���p��MlӻK�y	�j�2��d�o��EԋF��'b6�����y�\�pX�l���qe�)kHlѡ���G�o����U{U�D�<<zU0L�7�ߣe*�,��4snD�g�*׏�Ě� ���C�i���F.�+�,�{n���T�w�'�E��[�X�E��Y&���F�AK$*��#u���X���~"�����PbN+l���S=��ĝR�p���,��!�O7p@�\u)��<��u�MW��{���.�\C\��O�B*�%�����3�k�Е\6�hV`m�ilU,�Ma����ȓvM�6�o��Z(��g1����|u�rR�ñ�8��+S��VVSN���%��Q��ҔQZŘ�Y���G�!f5u�"������E=ϟ���/5����	���8R}�;�I���߬^X����wx����:�Xt}���Xt��o���˫�z��G�e�Ҳ�q��3 �{�����bD	�4��zfjo��n�b������J'��3�ݴS����B�ΤǬO@�G�JTʀ�K%5�a�UR��J>_[��0��Wu`��J��C]əl��!���\�C�S���j��n�F�4��f~W�zR�$==3q�X(�]��ѐ�b�D$�ϐ�9�i�$]�bl��Y�"�̀.$����e�F��j�J�w)�.�����ԹP�@�����"�o$��e��@���!��D[[�������!N2��
ǝ́TI��� �.sƌ�O��C���.�]H��]r��6]H���m�bz��p��*��+OooS9���'s��<d,�������Έ��=�^�`�\����#QIh�%`ҵ�x���
�1�'�o�CQ�/K�'���>�ޮxmI�1���R�&�pP5!4��d'b ���p2vT8���^tfm^R�P�}��PnN���p�N��0�G�!�c�U۸��ѥ�U�V�4��e$�۔�$W��6M�^�0�>��@t��
A��l���\Z9*��v�#\����(�h�a��0������-!���J��~>u�����Fط��Z�F�	��
>��6�V8 ��ձc)l���h�_��'�}��1��,�W$���3[���T����p_"���:����x���(;������\��r�F�MKeF�,���t�Q�K.Ռ(��;6������&������a(xWNe{�|M�\/w�< �G��$0�P�:�Yz��}��D�X�Q?���r��Ui\�S1��C�፪�T���Fu!�R�P΅?Xiq�䛚�.��{S*W�>��{ux-�������z��%�����ɧ3��k��%��^��a�÷V?)�������rr��	��Q������r�23�)�RL� f*V�̱�N�ea�X��D����E�ۜ�����sQ__뙛��필�#�CO����9�#��!P�j]o%����u`�EKJ��П��O����Z�v�S���j����c������Y1��Z�`�&��"����՜����sqZ�>�&��^b*�ov��b�9c�x��X~K:�ߒ��K�e>]/�ۚ�'���8������ ���׼�8tb����L6�Gś��0��6��L,a��\ۃF3X����� C�H%%��m|-`p��e��mv�h��ߑ��-V��-,�ng-<_5Ӽe�7�%N��~���MO��v>L�z��`�އZ^�s����o��"�k��(���i �BۙI�Y�rҝ��{��m���nGY������4�&�$���������y������H)���F�0l�$��K����Ћڹ������ ��w@K��#R?"�����}�=�t?�F���D�L�d��:�9ؐ����o?	^dJD�txL�b��8���Į��I�祦�?��������x7
�s��W��l��G�砃����m���N�ޕ���a�e��`Zͨ��A�4/��qW��z~������B�\i��{Z�թվ�̦�̼��jf��g �����]��+j�{d�[=���N�P���V�(��@(�/e��b��M�������34�.��=�<�K�2f��M��dw�Z��^o���w���uΛ���+�����慱ن7j�R󲘮I�x�E�a�c
6�Y�x&F��/z�^�{A�yXTG�����C��EF��i7�cS��Iދ��˭����*�ײo�������٘��~@�������Q^xoӚ,��>l�r{������B�����9�a�=��5�弢&'��.�_���������Q�V����_D��p�QYڴ�����^�6QU!�TB��J��Z3R`�����:ZH�"����m��� dYIE����'(��H(W ���4�F�Z�h5WN|Aq%$440�Ɏj�vg◻_i�\�q�'P���j�i_����m�q-=+k��y����9��k���{_�n��}ϠqY7ZcK��6���/����(�*L/���$:�|F\��7y����4o�gj��O��b�I����ϓ���'�6ד;1֮�Q1�O�	O�������<���Y��a������oo����{�0
ې�bywv�� 5P4�O����Ymp��2�:#Z�g֬��Q�s�2�D�Bzq	�����4�-U�� 3�T�?�ւ���Kɏ���g߻�	GL�o_��2h�.��*(U���o���ǉE�_x���Bl�I `��vG�@�A��zZM��s'^�����浺�������:��܀����en$q���?�<��WӾ�Xt>�ڍ���l��ku!���۷~���' &Ѽ6R�*�� �]jr�Jg��۸�YY�>;�$!�ug���o�tK�*V4)CQ��P#=��%�O���_B��>{�n�;�D�|���Xrǀ�!���Z2)a�{�a\�w�ߞN�鯾, �-��X��S�q������ż��eYN��<'��:��HMr�p$���)�'��s��`�-��=��2
�L�y�w"^;��U�K9��յy�������:쿗�>>s4�����=�P��2e-���M����"��6E�M�0,AQ*���;��ʏ ���U����(��Ql^�ǰ���9�!�2�Z�O��DM��1�#�H2ފD�7�X��sF��Y�\᥂�v�L)}$c� �J�7r-���wI��0L#�8DI)��)D�����A6٘�%�Y3z����|^VN:�:�'@K�SiU+��1O���n�-�iwf�Ra��@֝=��x[�"a���n� �����m�5��^� �r�T���>g�( o�x��<?~e�};��w�T<
��C~\+��\,���<W��k,a�k.��[WYD���|㍧H��Χ�+�+�V4�7^q�O5@�d`ۻ��#��=:��Cu)A��e}�%����ǜ�.��M��c��b`��z�FDS�ۣ�Vz���I���$���$�|�����}��Ro����j�Vx�wh�}�F�Еk�W�Ŀ��xJ`b?�C�^V����.�����)f��&�����?x���$��\�l�4����� 㤉*l~��A��9�`�s�� ��79��R�i[�m�2d��)J��q��s��Q_�@_�s�1���@ɐSk���ڶz(|;g����"m���w:��=zE�~�!�A���6�-���4�7U��I]��%�7Ze�"��]xn����g�v���:I�=��zdL�׷ɝ����Ο4���=2{� *�L�;���d�`�Q�"�t�M7o5x�5nhݕ-O�d���C�K�9`N��E�,B�D�LS�l���I��fD�M�o�ӱ�@k@a�|��9���~�T�_�!�}�4jDU=AFF1I�ߗ��ة���`�cR��+�w�JO6�jxT�x� yۊ��꡸��N�|ZQY+V� Zg�ѥ���f͂Y�'��]aЈ��\w�uU!��>���[�x�0Z;t�譮 ,���ό��?G��y$���2�^4�X6e��:A)�DQ�jt'�s:�&Uj2��5+��]�N���uBqpr�����S��dWM�|��o��=`��6��c�孲�r�2�Nq`ܲ<�3�G�_5��<TA�~(�|�o�@�"��\��c*V"Ϩ�$.0�AZ"�)�K�A�c�	e��7%f�o�H��w����V�2���b��%��-7�Vۙ���9�_�s�˭3]m*�����T�+׈l��m�B�������p�P�S��x�l���sg�d�=)�6��6j���\�Kʥ��L@'����]�j� ���w�帰������x�#]pӏ��(���>�oC&���F��tl�U�|��h֕�G��D��Mm�7(x*�в0]O��f<T�{�Ydy$����*�qD�����}L�?>�aV5X�!���`��i.Ӧ�2LP�C�	1��\��2XU�R2�����7�o��D}o��R��B8����k2L������P�C���aS0�@YbXu�ÜΫu`�#�^k�>$2@x-��F�̰J�ɑ�H,���uj��sӝ�&h�����ŏ΋UdQ��P�����.��I;绱�2�V��eL ݻi8)0v�e�j4��s�L� ����$���^	�r�0�E���2�o__U�(Gg�������q}�#Yqt��Y�ȵ)�$����(j.K>+x��b����T=8
�ԇ��`.)��T�����;%��N�5�͆��f�7�n��N�]n�'ur)L�Z��/�Te�<?��)��?���;OOx���,��S_l�}����JV��^j(Q��3��ݜ8 ��n�:�n�>��][��W6��H�EV16]����6�l|�Z�7��X�ށ��$n
>�u^5-�79��1�-�qH� ��;uj@�8,��aB�b�|i�c�e�]V�6z@�Hb|�w�����/�u5ϒǳ��ɝ���=!�>D���l�+;�j��CyF�m����Qk�TV�!GI.��|�o�n�>���p��F;m�5��ffC$^����
*����"�]H��q���"����0���e`,� �ֆX�]j�2�(�\���)t�����fd\���SCn��*L5�g�z�Z�lj���h,����+���[Ќ�c���MSrs���%���~����#��a�e�&y><t�Yt�n#����U��u&K���f�W7L�&��.A��$�����m�=�����N'H�ֳX�O�Jܙiz<2�%%2�ފ4�$����`VY7�����O4^(�3����by0�p�`.��maa���F������v��G��Kq�M��t�/�N��ٷ�U��K�(z5e�|V��.�ȣ�	�Kin�K��v�.7�qgm��+���P���%#�d�<r�ˀ��L	�U����39[�p�E��
5 ����-/����6��i�1��>r�z���H՛ĪJ�A^�J^�� k\Hԓ�[-,��1g��Z���^8�$��;����]���߿��`�����D��c��aڶn�t�IS�u�b�;���|+��<$e�+�m͐V����dc�1����y���W��Y�4�=��v�f��u�T�4VA��F�&5��>����M�>(��W,Ȟ"�*���1ٰ����MYN�Z�OֳT>���w*iQ��J���r_����:�䬞֥e�/�!�f�'{���%��
C�kL�m�� �6���:Dn�Y&C��}���q�T�a��#�Z0z<I������1fx7���+�2��D���ȨH������7�?���9X?�����v鈌2�/��x���?6�jw��u���F�����G�3�@t!��"�1V&z~ڨjJ����ʜ��&��r�2\�L�	8R��a�e���q�1ʣ7�V4���@�cto��:�뎿�����k�B
D�%\p�+�h�	�\�7R���X�>�]?Z$JT��D�d���|/ނf�I���eYLy��"J��CYSu� ��d�� ����O�Y���o�ST?� 8T��tvI��[L��݇I�X��oMٛ�B�"O6LH9����)����ޑS��)hzq�zV�؅���FR��ѹ+�@�Y	��GI�v}���+�O�U���k��2�޵nk϶o4P�,��;�5L�Z`�|+_)�܈�[�l���,<��:=I��_�	yd�ԓ2�m�����w�>/q���%l����T��8��y�U���~��<��t���b*�[K�Dx������N �+9�a/J9rS3Q���x�� �l��y�kxҘnx^X��(
�c0vV�z+�Ȝ�8��RL��؏f�T)�/�>�dOLaP��1o�N��,j �l�q�0So��x�5L�Uz��1�X��Vd���i��q�N8�7+�Fd i��*Yx��BGY/�->9��3����ߜ;`� ��J��P�ώ�kZ�,��(�x4?������^�JJo�x����/�����Vݰ� ��vuO��;˭!�$
ƻ`�����	�jW\0�h#��c��ͷ�?��J x`E *$D�u.�~!�ɓ�? @�)`(vD�����o������rG���
*g��H���N�d*1��Iny���/BD"��l3�B|�W0�y�5/-��=�T�&�������\˦�� ��sh_KS���H<˿�<n&����(桾z��P;"I�5���V��M�nK�-��羓
�寐IROԭ��#�2�B��]����*0��T���kb4Q�oi	�'�٣�f�@�W��ܕ$ֽ-�_�p$�I���`BF,|2M�I�(��ѕ1\��k8(ٙ*�C.�/�Ucf̿��Z�R��P姩�F�Pq����h�6ߕvM�Gј)��$��Z�j C�8gh���^�U��i�U�p���� ļ�Eh�'B��y������_�G��@^95���`L*:�Mp�NE=<�_RϚ0K	���9C�m�M����@�HÓy��b��!�PIk�	�WDe���<��eH�"�iV1�
�YIi��B���ޑPCxl3�AM���  @ IDAT@�i���Ӫ
������I�Sح"��o����]��WOe��,��ƸO�"ʨ�oG��=TM�$�l��̺�� D'Zv�-�e�6ΰ� �c���.u\IT*�"b-�ƨ��& d#ͺr�\$�y
}PMR�89=�
"J��J���Oٙ��"x��v�q-����QD�ց���� "��/�/"���Fn�ԍ�"ɪËs���Q`2$�!�:y%�(��%'}��83�v�����D��
s���Ttf���$d^L�%�ץN)HND�ԃ
'�j�>��:sd��4���8i����㠝���t��&X�1����:\˴0D�@�ȁ�������0��wFK'�D�"R����-�"I�L���*|P�1�%p:��;�N�����2�.,w�Aq4��j�������C�|	�=<��D"X�K����*��D&~R��e$��Q�����L)��ȇ��^�0�`<���B&&UEɧ_H�?�G� �{T��<��%7��l_��lW�T^����PqU�R����2P���QQ��ƋqsS+W�dQ4!�@@Z�8��7�*Br1%���N��I�h�W��@�VpT�"�&6��b�u�}��Ĝ�RQ{���=������*7׸��!�;�E��J�jv����|�	h��Ǯ��N+��a�� i����ۻ��dab$�߁[fi��^�'߉��j��a�����Q��&��-��{�������p���� &��o+2{xTE�v:�g��+fJ�L�)\cC��X��C=O"9�o�g�'6{�6��Q$�HRKV"N��O���Ѽ��)���"QIZk�ETBD�;E񮜉^@(�+�$d�����g�����4��_�X@�������Z���W�Э"�[@k�az_Ք�S��� mT� ��?gR�	���o�	.���w��%���/�JFi0bѪ'	'e����D�7Sqmȟ�|�ԧ9�Uy}1~�.��s��F������_�+?�����|���o*�w���B4����w�I���.��kE`(Ơ��Xw��;f�:�,�+�I��L��\׼�E�J��s�p�j5�64�$��&�`��Q��]X�(�(����r0k��*D�����t�. �B�Bu��#�[��.%�_� E8̢�84YB�~����er%	A���	F�g4�7	A}JH$��=��#7{�E����tK����xI��
�
��V��!b�=�@��Z�3@j	�S�Ҙn-{P0�� "�A��"JEXa�0n+":1�~=�O�y;�/Z��q�(��K=Nط5r�/x0����q�&]Q�wpK�7�P�� ���R��|���?��?�`�n�IPI�����(� Ѡ��Q۵i����eQ��]9o3��2;.�!J�YH.TNq侄Do���!���ϋ��]�b��;M�$�FI�ca��$�H�;CD��0:�jIH��Ɵ�T��J(�i���\7��g�h�.$L�-�.B�s����M�����:�_>
1���Y���U��)`���@3>�|����~��E���o���c� W�4% R����Ԫԭ����|���`x���.��U��8<oh+���htF��Js� ��>�>�?a	B�_!l��$Ԣ����@]C)�"#bb��M`nn"���h#�B�˛���u��։���3�CL�q8#P�=�������N�@/�Q�T����Kv�ς���"iԁ���������( ���'6�'q-=-��=�[m��	ӕ�\'BkI/J�!�K��p� C�U��W'SH{�ڴ/5\����1 ��7Ο8y(e'�a��Y�\����E�F��V�D ꧘�3*�C�:~��ؾMc�!LSu̉��0�p��w��G�)��-���$�f		���H��%`�	V:T����&݌!c
��o��;��;n�Q�ȍ^���PtW��y��
��M_}WӎC!b�oR������ED�e1Ⱦ�.ѿE�ɸ�e�#��`�$�7R��	���$$,V�(LNI����B�`�H��t~�KLy������&�u,����v���sk�Q���1�f$��h�I�!�@-�9N0���I�qj;tvH��u�Q�ҶDNNC��� "WH�Q�y$�%D�Y�`(���p�ix�L����i��������K�|K�@B���*-oh�����5�O}�,�"�8U'�w���{�����G���P/r�X_U�v��E�	V��+�����z�o���M��/���s�7��i��k!\��-��-�n�(Qc�Z�M5����2+]�j�/n��[��w��;�%�g��]8�5�I(#���#*��!>��L!�� IVI���*�ރ���y��ZDN�<8����pC��ɰ/��$�$����
1YC ��u���)��5��tQ=6	e�C|��A__�]����[� ƪ��g�Z��ʄ�H+H���o���+�E�-&��R<�4m����o��RD��_˃�s3_���,�"Nmo���F2��	1`Z��5z�i
�v�*��Tiv*�ꗊ�=�ρ���U��^i[aѳ��.sЯ}A[7�e���ջƛd_��	���E-�>�[8+��f;���D�F��:�b�<�ב ��� ��C�r�s"?>rW������L�+���^��^�S<(�+ j���TX���������	�EZ*Kr�[$5�
������We��U:uIn������[�yU7�RR��ߪ��y���H� �d*�{`c�.���1P}B��0�p�O����Bg B$��j�Ø�ί8���1���"8!،�>+,7�� $ ��.����J���R��#8+X�|�nO?���o4�K�yZ�f��^Q" �ZNu��O�7���]�5b/d��4jp�hD6��B�S݌�y��-@��ϛn�+��w�j~������������+�h��6^��NkUT��:u�	8��z�ϭc����q��C�����	a/8�喏�%W���3j}G��u$:�wU���!#�����n�D�埯U���Z��#m	:��b�ጄ0w���ZqO��s8d <�:1�8|Y	��k�!�F�q<D��'B����w_��}�Ѩ�W��Ec�I�@��\�ϤSS�!x�ꓔ"��{>S'��{JgN�o�R�ԣz�]}p������.�9�;��5|�B���AڍS��y�/��jCZ�#L0Ʊ�KZ�׽]`�ȇ����?�T�������<�-�S��ŗ؄�n�[����Ru	�Ka�e��<L0�8!ފXl��郛V�H0�K������
c�o.���1�LB?;�i.�'蘮R��J�		��~��mzVE�Snܫ/�qc���; x��ޣ�]�	����=�#͍�Vg��1�9h��]/�����Ox����r��y��и�o�ܛ��?�n�p��b�ј�p���[+�Ol�Xz�
l&��[��l"���e�˳�%��Os.��v�&�ȴ�^�(ь%������6m�$!=|��H�]Y��[%��5� ��+t9�B�B�#He	�'+K���<I|d"m#љ�,[�5��/��sPH͖�C�S䛜[:��M���IZ)���&��s|�(|��.	�$�[c����ZM���vC6���-�$�\H���rp&�K̠E8�bF�F���*I�D;�	�)�Zp��E��P��Ӟ}؆��������Y46W�WH�ʙ�Wm||֢��0p�'���}�3�Y[�w�c�xȪk��+���ٔ�8B��lhf�H��X��2�TZ^�ph�� ��Cu�����4%is�CY��*��D؁�����&�K��z&4�|�T!%h%�g�)S�cQ�����W˱�6�	�3]ￋX)o6��u���Q��O�a���������G0*ͭpZ8%O�YAc���B��W5^�x+4\LX��F�����@ӄՆZ�����r��ς�����yl:h��K�vOY"�/ݯg%Е�$eN	��b�H��bMw�\9)�������|��y�j�*��;{
�����_�4�D�O|�J�OYv9W�u���-�ɻXY��6�r<���ϽlKs笓��ο~�^>v�6o��}�,����^��sQ$`�H�z]ف�!�bxy71XuZ��`��E ��� ^�$����v1C��K6R�W-���ϲ4ŤF9�A;�F*�8M��i��	���&>ޣ'5� 9�� d�j�5kTV�����HWVHL�y��!sA��5ɩ� �[����1���U#AL�����0�>�ȱ]��(/.���i��;�gh��)9tK!%k�/PW�J�M&k6�iC�d)e������n���Gl$K�	��9�d7)�E�bGi��j�_z�ڜ�e#X�]�ª8���r�Z��-^|�|�}`�|vh�,G$S!��~v4����Z���/i!��SCۡ�-Z�y���06m_#��$D�(뤎 ɱ��V�:�E"8�yͰ9M&��A�&��1 ���,0� ��~�X 1��~>�4فIM�����bNb2�����]�D���6�W�m�_���_e��k�_���z]}������p��/�v�h!$�7EaЪQLG�NᷟY+��}�����֙�E]Z��5m9�7�z0�x(F!�ĺ�Hr�MM�$�QZ�h'�ll��v<�@�X������S/�������5����~]��������%R����[ߴ��oXy� ��,1�����B�@�?�6����:=bY��-]<��A��9�.��5m1[�my�dG����{���%Ӓ���P&����$��a0�@���3PI9e/u�b���
 ��$5b���@�aa��JΖb�!�|g$�d��!:ܴ� �lr�vr�L.��!��'3PFZ }���.2qH�:Ie��&��8	_j��#���g�nMM\oc��`��Y�� J�wH��+��I
۩e�̹dU���b���G8RPbh|�FI:3�Ve���!��q��������K�N����΂}���Ƕڎ(�F4���=��#�'�۵+' �椨a���њ��fH��!"׮T�\�����%��`�	����j��6���b�h�'i����",���O�kj�47q��pAT�&����y!Ƣ��"�Pj�RP����>��hFRݗj�A��	�{d�{Mcp��[����	�������m�Y��5�X�F�{���oO_�����4\	#��Pq(���n��:�TqD�r ��v�h�R&��~��C�tt�o���A���Y��%��yE��,��P�j�%ߴ�s-�V�j�]��q[�W`�l,�����N�v��g���O9����V�U~C������'��3�%��AԬ���)�����n���!6��
��f���&��m����-�ذC"�Tn��_��s�l�cԗ6VI�B
��v+����s�e�C�I:��=r4CZu-1Z���Ц�mI�7� F��b⠢w����LG�}D�
q���N�ԄOR�l��� ȍ*��s#�n!��w�Q�����,�c��$d��
�,Ӣm�"��Ҙ�ǘh�h����a��sf�&�ɓȄwvO��dnp�Xb�B|E߁�y$X!˲%�8ޯ��ơ>U��@� !��G�U��g�ɋA�|�r�c�Yڰ�)�%�py�dW�V��?��r�Svy��'�)��x�35�H[G�D0
�4#�Y`�B(1,%��`�/Kcz��mV���1P�-�(u5�q2��w�����D�����V��P��	l�0%��"m�9�jGhV�E��:��J�]Nr71a�~/�F�
p7�oz�Ϻ�gn+\���_��L����nE�F�|�$��P�U�)u1��:E�~?I;���C��L��I���hMb\|���6!��eU9�eb��h��j�)���� ��o=�U;]�D�T����D���K����0jR�gL���E=�ڧ
�Y�[s���O�]��{e�_��'a�Ǭ�o�ٹ�������]�����]�߰�$�#	
�@]v��Hٵ���)���T��-���k�׬�T�1�������ՋgN��Ex�~+,��rL2�yTYi�	$30=E�@Eg� �L�;�7�i�F/y��5����	�3P���� �`��@[оҶ����RH�L��� �`�.I=��Wʵz�#���u�
�gΊ@
��gA�:�QZڋI�"JN�|�D���I/�2풘�	frZ����plO��%e&�������rpR2&ߔ� ~ԙc���M�0ш`��*}�]���u���� Z���Ǣ���P��R0f�~3hne�Ik����d`\	:u�WpU�a��aO��*��xh-���:4���q֤@�p��A�8H�;�U||5m'J��4�<C}NH�+5]K����-BR��_��x� �5}#��S��ȟ����y�mE����}��q��,�����w�G2�a��XE�<���\LME��SEL����i��X��(bF`.�\���46���wh ���'Lf�j��^&! �~�)�����*BB���_w�3_2��O�	d�����4�{n�'.d�pèm\|_e��-\<fo�>��LҌag�9��羭$8�Pa�Dޥd��@�Iqq��>u�^�^e��4��ڽ�l��ɢ��vܥ3v��e��{�I�$�6�i<o�5�`���}O�e��Q˫D��;��65ƀ �[^���*�OH��@�1 ��˒=�R�4q�v]�
�D��[�}[���t��DP�{8�I��@U���|X2O��5LL��ƥPo*&�+�0C���� �i��9�bҫ���r�����ٳ"&�z42=kd���p.�����l��X�c�lr�����w[L�#��i+��.<�;dl�'9�,p��0��ux-�n��͖D;�A׉�m�|�cS�	�S v��0.�Xm�)%&As����i�l���|1�b��J��p�����3rJ���hG�J��4��96����w���d���ۉ�:DP\�~���ĵ4 �"o���߸_�F	>�8�Z@��(��~�����祭�H;k�X���b��������2=�����I�,hD����;�A�P��=��(	�t� <�G~8j�C�2�I��F �M�-�ʐ�4�B�9�@$�ј��d1a705�� ����;��1�[k�Gګ��=,^{�#��h��"�i	a�TAAC�!�$��o�D�B�VB���C�4���$i��W�dIn��_?��I؎=��ҕk��RL�I�j����q̎1�
��J���c~ kK�Ri@�)$m��A��qܜl�Z�����)CU:�k��(%"�@�bn:�E *��q-C�e�qoEcSu�nw
�ޕqR�A!v#�B�+Suk�FүKJM/n;�a�[�x�4�#�k�V$|��`�$#.�-�qL�1�����[�9H��P2��],���rކ��l�4~��i۸�,Y�lrT�
���>0�*�I�c
��s�A�Ƞ�u�����%�d�W1��B�k+'g�,�B8��(:Pv��HIꮾ3<g�m$�"A�hW�a�Ⱦ*b�Ӯ"�����db�Zw�?]�nR�mi�G$����d���l0AEZI���n��?����H��h�����p�0}�A}�D��7�~J�SC��Ie���d��1	IwZ�ݟ�\�W�m�I���3��o_ߥ����K_BP<X+!A�c�>1~��/n��i-���Hr���ݛ=��\w~Y{���*�[�h6�dsi6)�)R���2�E��G������?�#?��L˒b$Q�D�$�dod�X����
��˟�7o��j��Iq&�[���޼�'O�s��ɓ'�&�(Dp�)ޡ,.�q�l�,�|ڜ�N+ծW�"�&���_"��>9����X<��t�Vf	���?Y>�������7����b�dYo�wt�1A�U�?j�a�ģ���B�\,�s ����Q>��G��'���ES:�q��;/�����`Z�<Z����b(4zp�V`f]A#Pp��+\u��O*FX������������FY6H�[0��)�+�-�(0-��K��2��J9W_��<�9w<փ[�֝�0�a�2�
���24��L>V��Q���!8�4GN�:���Yk
!��<�e��b�9��`/#<V.�ʁ $:���O4��ğT�Bh��LF�V;H�F��pIS��2Y"v3�[���	��*h!�q����̬D��	�C	u���!�i���j���$�:6�'u�.B�r�F�0��M��[�b[Fp�S��kP��ft�V�&�n��[aN��{20���A�ʙ!g@���2}�qg�Ng�E�1 ��iW[ʴ�5���1w��$'0�G� 	�
�wC�k�Q��&C�`���A-�	�@��8~x�6rq<� |O��ރ�#(���g��L~dj����Ƀ�Ɲ�d�?D7e@��ౄa�r�AJ[��������Y\�͉Cׯ�K�n����G��7Ε�U&��6�92��22b���>4< \Fіp��u:t������>�k.G�����8�5����GOÂG<%(ꍝ9����e-�D�j�Xp8��ٖ��Hꬿ�����"؈T��R�������ЀjZ:��j�P�ߩ�z1�:"�y�;�?��L����wa�^JO��?EU��[E7�F�u#�� ���I�o�0�gL������|������??Qv��������3���r|Mbh]�8|�UH	S�*�8��Tn��ih����G�]��M
s�Ñ�w�G�̎`aJ� ����W�����  TFT��H����U8�ޯI- H�O��v�p�J�L z����
� $O��7��֝�)�B���.7~e<ҟ]�1�/��3�w(H[_�I��Z����j�S���M_�Q�L���h\�'��A�rī�h>�N��"YF��{��< �Ux8U��J��	�ԃ.	90�r<z��yH����ߕW^*��C'�u� ��p�à=	�9Z�h�@�r�|�`d߶}4�s�,�=���e|{������$b*/ ] ���w�a�FEԐJG��;2���:3�P�m��Q���]��z�?�����c�#8�Y���dG�^�����Te0�#��kE|���Τ^�{uL��)�w�I�~Z-a@j�D���<Z��4ׁ��:^��()6����;�4��M�>�O����1P�4�zƿ�2%�0�L-���X�KU� #��Q�FY�
 ��-���j��b����Vŕ�UoMJ;~�y�KGvA�j�<���18�U���<���`in���-���6��&�E��k�
E�g���.L�!�Nc��ٙB9h	C�����S5c4E��'Ki�D}N�W�S%`�+��\+�_j,4�{<�f�_�7�4y����<��v_�k��"�P�N�{��v�g~w���v3�k�@�HZ��ɶO�)�����{�T�u�1V�
b����Ҳ���P��W��͔�׉�����!�
=˹��r\�d�<ĩW�PS��\��[�PA?��2T�$�<���ż�{����f ˹1�/!��3��V�1�D�;��@Z�A�eU���T5��,p��ʎLgwp��{"�	0Ƒ��V��2{q#|x�ۭC$䳣�t�G�6�pe�zG3x��Ǟx���2���"��vO�.�4�x������x6J��A�u^c�M�!��Q���7ik�ph9WmԔ��:2�X�!�Cl�My1$�]�Pz BW�QxT��L�Z�ݬ��F���A~��M�.��Z
�,[f���Y��C�o��*�D���"����m��DY>��I��"��@�@ �tC[]�F��PYz�+��!�_�+�,#4"��//x����G���!
f�w���+�#ީ=S>{�Bg�
<Pp��)��b`Y����rjv�j�sx��ҧ?]��o_+��qvKn�j��8H�em���$�cxm��Na�<Q���9�0�L�D�Q�q�A$,�@�h�B���r8�E��)}G��Iw�O32|��u�Dd��󧏃T%4?h����v �gNh���{�>�W%n>�7@|�v��u�FX��H�v��G�){��NRc��c��kWkO-�b��B˼���F8F�#�7�{�C�=�j��ī�҅�e��?Y6u	Xa�����}���P������m�R��x��Q�W j�?]{+�0Y��s�"�2JG��F�%|��á<uDL�����$�A##q�V��#�:0x^�J��ıK��L�2%B9�UW}��#�3��oK?��o_t��>daH�Y����n@��Wa�a��������Y���8����mZ�G �w,?:tJa�Yz6tF]���o�
h���rEw�`�[����q��k?�:͐^��W�2���s������ w����_<����|�OX����Z��W	W��F�������'p�7ʣ�-?V^\:���h�>1�ނa�
��ɍ��:�I�Q:��OP�_	L�:$�y�7�r�5�"'B���+Ԁ1�����ewe�S��r,��`�Ј�<�O�o��'GY��a�$�CB�Yy`v>�\�LEUx�Y��.�����X@������z���໨���'�|�ܸ���ֱa�l�W�0&;g�.�D����a0����dF���!<����6�$'	�Ĩ*ޒ��a����34�{X����	�;��l%��6����N��aW�/���1y�����E�Dn^�H��g�~�v�$a��*$k;�mRB�
)1��;�q3�w��q���h�\;�v80P��c�J�{`�����i#}!�H�>�I�e���˩JŢm�O�Ͻ�T���"��aʍV��L��+�5�R�[��i��@�h�!2N�B�,ød7ő���~�< ��	-�HB4V�0��`��2^�3W�s/<������-�.ymj�z���]r��U*�M��~��[�,�<)�͓�iC�!EDW��)�v�Ҵ���|���o�?Q�cv�i����>������ �?OG|�c��ꈲj��ik��g;�z��ЭY��=�AA��&;�/���8�̞�8�a�\ue�~4��XGU^�,=5]-��e�oWX�� Ҍ����"5��֜c�g����8��'݄	�:jY2��gl���4�!8D�.��5Ĺ����r�G����Q�
ō�&����.R�E����c�#2Q�7��|�j)#���7u�4Xx�v�e
I���
�m�t�L��+&
�b�1C2`Qǚ޶�A����|�!b�jS~�$����_"��T��z�窘<�r)O�	� \�nV���j�2�=�l���M�����+X�Y�rPgD��첒�ȝ3{˿����:�N͍S�����!6���dǯ�E9��Se������`��^-�s�������@3�s��l@��,��1�'�F	9H�O�L����j^�_��� V�w�4ɲD�)���C������?�7|�]9�l�������W�*�~�f>a�}��	�ާ� �%��6�27str��ۃs�!���{�~|&�c��l��6]�����C��h[b�N��D������$J����o��0o�f��PU���.yy���;���#����Jk%�"����F� 8+J!`S��%t�Q^�}˓.ү���K�BkN5�9*�a�`��_�D��ҕ9���i\����$�Z�ck���c0ꔾ�C�d�W��ϻ%�@:܈jN�9��oC�b��:�'������w]�m��c�k|�f���Ă5�F�fOu>�[��o�[p@}��<>�y ~��a�z�'��A���r��y�K�O|X�x^XgTB�)�Q	�����Tsss!hm����X�g3ނ����������H,UB�P�����`�[�!�j��;���l"�g��+��e`���;�5�ʰf�j�W�T�����[����4��+S"���Vc`�=XL�P���xf��=|��%*���w�
����6��`�ă�uJ#������1�}B���d�v{A��8'U�-3���Xa�����>�xܸ���i~���\��_>q��-��8pd;;x���a(�K�.�����O�9�,�,u�c�AS�Ne�
�l��h�����&1�ٜvXN.�����+�.�}���ԏ�P��lW���2񏑩��4��Z/���
e�;)ŀ[��Y��]�\W�$X��B��OlD�Uu�w���}ܣ�����*�zF2`��7pR?uF��g�����CŁ��<xs϶��C��R���I�Z��4Z�N��q�~��[����D��p^�I��U;�ܸZ<�0���$ӋQv���o}�]_h'�4#�p�\���e�y�� ����<@U��;��������� �J7�c���P�~ �pԏv�~V���S��ܮ7��Χ��Aj�i�w>���(�<=��I�e)��˯�/�wkW���?�����pJ�g@�����kȤ�+/���d��vjp��tE�7�NI ����f/癙��W�Jڄ�"�����
!A�tp��z�u~��!�Fى��fu����j��M6^�W���⬎v�
P����b��a\���L��z�.��J2���@�¥q�$CeeC��\U@򶈡ٷ����0�:\��S�\i>[�ɛi��,��S*�XR����Ee��)�N���7ae�S��<b%8ֈ\J-ٲ3)lU��R������@�0lh�	_V�(Ȥ�Wa�T�/i�8xh���˫ qӦ���̥2�7��.+�Xل��d<��1���?p�\�p���Rå�U@eƷO�PDfj�����M-�R���n�S:���r;*�n���VW0�����ޖ�U�{����*�����kg��d	OR��E��{�s�^�њ�!��D�����l`����; Ѓ/1�Nځ�Ɔ� �Z�i����C�%��#�����u�u#xW�r�
RYW���YA"�_G�ƌ��],S�̡;�6�L=`��-��Z5�\�^���"�g��F�n�W�P��Z�k�D� {�ɔ	��A`��[�!�5E˴d��3>���O5 ���}.^���Z���x��qZc���W���mt޵��w��h�J}9���N�n�Q%�;��v�oq*LN�����.���3���iXҪ��6�ml�ڻg��V<��Ү�I��� ���%.�h`b
\^~��E�uz�DU۪�P���2)5{�b+JC߻%�v�)��^��]�-�{��3A/'_?Wn`����j:t�>V38��B�4ğ`�0�W�@Ha���=�n�D9�I����x�	J�
Æ	jٕ+���)7�n漐���K�K��X�7��G
�*D�b��^�Э���2ڒekdՖ ;�)��
4�I�yԄ�?LHz�aV ]rz�����PxȘ���5xW�e]��z���;x"���y��[ۭ���mp��`��'`��=�~�iJ!�-��,��BE���VG �1xm�XH����(�Ha�Y����o;��C��)[By�:Fѹz����LM�>6T�� Z��.R-���=��x*�74Z2�P�0���!	�`���\Cnj��{"򭒄���/	�*{V;����7;���gG���Iݨc�����^���Zkg�0������r�Ӗ�8�p�8����9º����>������C��=l�!�:����@��Q�_r�O�9;t_�k0g�}�|���3�W�����g�;3VoȊ[� ]ui��*�1;�J�%J�@/� t�����Q��@=��$��2ݨD^�-�]N���w�l\�Q4SYH6���i�pJ�F��+d8!t&��^�0���k5��V�j�d\��^�����I�xjCi���+=f�u�����ܶ��Gʬp���DB�/��y4���;j��ئ�>7�Ң^��t۹��FHH���l��D��ݸQ����|$p�R�Cd�س�U[5�����j������D��=�:wA�����S��`�C����R$��B���?�
�b���*���x�w�7���溪e� ���	��a	l؃�\⬇�."<<���
���Y$�&���\���j񾂥�TG�,y��d�		�i�<S��t�⁗-S���B�y�s���4����Zߙí�¨�a�r���6ShZ��h(��t�A���Ru��3�Xc�e�{<�� ²�7�)K���0O���R3p���q(��U�d�BF�e���j�yE�`Ŷ�N��tmSXt`�em�V���A�m$A�
���DyQ�i)+���Y��|7P��ג�*�sf�;��������6�3���0AyU����~��KD�~��Wʇ�؛����m�r�k�r����o��c4 �o�*b�P�ٓ� ���o[�3_�E�〩���o���KG���\�M��?�9����]f���Y�z����~�ǌMm�����0�ꂊ$0	xR��!�8�8"�ͤ`	�ŅQ��-޵3x|V��r/ޭ��L�C����+)aJ�`>7�E0txpdt������2�Ϊ!;�z8�m�
\#{=�n���L����t&���Ա�F���k{`Я r��"�Ȣ6�e�#d�k��G&M�ްm;�y���02N`"Vslǐ�r3e��Zh,G1&�����T�6p+���P�(u��ԅj��{t��V��h��rvh�k[�
��>[�Z���<�H�M��\��P^;}��9���xQa&!����<����6�Fzw�1�$<���v��S��Ȧ9
@�)ɩb��I�-�^�vf�N�t�rG=l?���^�x�r߃{�Q�p_-0F#7�ON��J?O��s�/Ek�b�����C�G@�ai�]��џT����[�B����������ڇ��͊�~`����UԥR˩"�)�(ޗ�0��:�1�K{jBNSW8K�>vg(�ΧZ�K�,($�4B
�C�Ux�\��'�����l�J�@��TxBS
�0��܁�獖V��a��N^���7��P�\u��oa�?�fˆ��v�)����p�r��������S<�oX��L�f/��m�6)p�D~�#�ۀ�yZ�톺r�"��'C`��Q搷�UFw������	a6Rn̮`x�aNk��f.�^��Ʈ��ՎQ"�,3��&���KgB\��3��r�Èl&��\U�U��hXRm^�+�;v����Y���	b�S$an�`K�����NHUI�Y"ݹ��om��4�5���|���lO��z�Jo>���_EŃw2�t�נ��� 9E���7.<��`��2���I;VΝ�R�;Zv���Ybj�:D��12c��_?��F����e��t�Va0I�Ƶp�H�d�!xL">g�Y�@����u5��Yߧ�u�n�<ӏ�vzm�n�I�`�U���Ht
�yeh�p���P� @���8_!����5|J��;x1�˴��U1�\*��&�ʒ����¾J;$)EJ�F.Lr*���Ĥ �(�s԰0��{
��d=C�*Ux�^�0Z����eP%�H�ܪ-)�����9*��/ m�.��4�� T������F�H�؎��H"��	��2WF=&X�X��u���_�Bٻ{���'ĕW��n�N�����<۽
��")���`;��:R�_�x��ou�< ��*a�q�Z��n)Ҝ~*`����%6[9ۛg��$��νq�[D�����Z�ҧ��:g/�}4Es9��ӉZ�y+n�(G;Ȓ<~�_�#��]K�n쪴�u�	q��Q�}/Kv���s0�=���h4u�k"��ix�RG۪5��$}i�Շ"��ˀ��������&��9�@5�٬2e`�N�b0* G��;}ɮ�h���*����JrLW���. �'6¡�WsG����`�k�  @ IDATc^�.鲫I-B{���D�g���	�!�_��ǟO}^�joh��g~�^oV�
��Bb�\�����q��������2���"�6 h��y��>�#�&��<�"3����s���A+��y���A9x��R%���Ȭ��Ƙdh��o.c�N�H��������.o���w��ݲ�&	��ԣ�����K��5�X�9��C��3����1L^�y��9;�=�����ϑ�7g���BS]��!��������*�����*��8�����b�����q��X�J?��lC+#h2��>G�"|��*�R���E���A2���*���� ux�7f���N~��z�"9y�I9��
���DvG���Z���Ԕ��`����̺T&����8-�q�Y��zzX��J:i��kB��E��=� `�^���i��S����o]�a1��3´֙G}��ģ�Ƌ�׈S�����D�:x���n�:yj���	����j&�>Z�BE��tk�ܸ�^�p0���3�������ݤnmQ}M��-�!�wS�?Jފ�F_!:��	��ͩ�i��O���	C�����耹����s.s�4�X���A�x��(�>=����6�lC�#�TM���˿B� �/�-�9}r�������ahGw�4�2+$`>�Y�2+*uʲYObCX#�����N�n�^�ꍞT���A=an �q� s$����zP�)˩�4��$�ٺ�#�Wܖ��,��?��ܫ�⇆u���w�$�Y]�v7�^a �´�\S��S�zR`�^�U�Lh������B[�a,�
����:��+})L��mS�W�-U8Tbp�* F���Yl�nhEXd^�sf�,�Y��g0Tzb�bپ�e/�2Vf�Tg�3w�-W9���e"V�Ca��������.�`�"�y��Pc
���ɼ��_Q)�өXM��VM"�-R��婝PD����]�q�]�S�fS��qc�u�_ɦ	������:)�9m�qf&� ��{Mܥ�tOF��������_��-��wp��׭[�a���2��:��/!�-���bM��cawm	��h�v�C���˩k���m�Rf�����i��S��h��E�2>a�؎(Oo�%���Q��BG��tX�݀�!!�Q�C���Ԇ���:
�Ҿ�˺j`ݼ�ѧ�]f�h�~�1��Z?�R���ʻu�Ꮖ7�Gմ^����2z}�;I'�������/��y%�_?E{�mB����ݜç���g]�*X��7+5�h�!� Z�mЁ��\�6���vgϝ�t����@"F�ۜ�Ȫ�.>�B]�@}(v�(�?p?�S%�R�+������u��oy��u��ӟ��7����nDe��w�{�S���
K�l���v*�����6�@���P8.�hs+��w8�_�H�ec�e���>v��?eZ@�Y_u�{'���
 ��D���Z�W�T��&�mNO�Ԁ�$�u҄���F��Y��Ǯа����.hJpb��}*���h��S�8���@�T��m��̈́�,/6*� h��w2��kF�����7�)�vB��L��e�����*�sч��d��@tp��
	ڠ�4m�p��G��SkJ�j��K!���)�ls�]����"�9��D�Y��7����KNZB�S>q�݋�ѫZf=t6۽�f�γi�3;�D��oI[��٨-��S�D���^w�����������Zwը*�������:R��:�V�Qխ�V��:��(�)Ȉ����^�(�*�Z����]#�6scwj�����8�ܟ|F?�O�{�Ӑ���r���S�����\���T�� /�#��h�-qk���ܫ����;˯�"�v���Vx���/�?YF̚6q.�a�M�����ΉD&�)@�AJ�0*�LP�q�Z����}���7jR�dky�p/ +/B�j�Lf�m�r_����'���]�ep� Ȳ�-_��:�]��a��۽Wyú�w���C(��tݡ��T��>��T��6��]G�Q�a/�g?�+�W^)�����>NxS�\�<JB�/����q�#�7�3r�x���l^UW/G����H�V��?e��X�{��zs����O'�+(�ʱ?L�W%�J�vx��Ж����O>�owmޤ�`f�9ٮ�FQ	�e��(���V����iQ˳3�S�R���;~F`%o�����ٝ9�|
w)*"�|�@�l��°)H�@�u��2���	�QV�<~6���Z��i��������tʭ�V�iv��vi����.�ܼc^��ߜ���Y�uy�[p�ݖ���V��k�Q�u�tuD���%�FzK.��<]يb��؇�]����^C3��*9���,GA镕(q���&�����C,@��2ݤ1j�qܡ�ʳ?tG'.طX��ȶ!bEh��f�tb~?{U���I�#�Z
bZt��jh^E�D*�cEl��ag��TZ�u]Ѻ�&�:��܌�=���|�b[���ĝ��3���{�	7��ջ_o��������Y��l�W_���7 ��O�+/]*��?N��9mf�~6i��N�ab���sųD!v��S��z8��m�8����;Ũ��"�#�a:�
qa��V�m����K��7���( t�#G@�@Y�r����"��m�
����f]Ӧ�;(n��յ�5F��rH7��:����d���ܮp�v�k�U�D{�zꊀPP>}Reǣ���$�㻼��V�pI��O�i�M�t�>o}�m�&�#bS&��3
?F�]�噊�T!��]�|R5�Z;����n�.��՝7r�P�ɾ��q����vJ R<�h��=_��_�\y�y�u����������*��r�;jUJ�_��2*9=QU���"���$Q�-UB��û��ٽ0��g���8"5����Ɉ�d�	_�(��Ƴ�s؇n���ݸ�L�fZ!aݾ�}��:�9���:>1���ݶ�P�v��7���|��Bĕ	���h$���!^�j*���=�5�����<��|Y�6�bim ���f��6`����Hi��¡E�vDF&���T��K��2�����Љ|f�(m�~�nZ�����O�|ש7hI�N75�Z�]ʌFB~�X�%��nY\Ti�P��ju�NVG�,���o��SI��R-�\���i�j�F�_�a����3)�G�c���w�W^�/|�Ķ����Q|��R46�Ğ�!��>����MG��T��6���+����Z���$oZ�ȓ�?[5�;�[r�k6ӝj1h�Cl��}sX�hp��NG��H�6֧G!�`�?����J�x0,Z�N�Db��m�����I��X��95�)l������=��%l}a��~A���O�W�*Q����p��	]��4b;Bj���,!3}JI��,�|)�g�����p[G%���>n�A���MRQ}��b��u�hpj;S�+3.��� �2%�@5���:�g~tn�=�\5���(e����& @��iChdL}�)^I��w�Z�;xj����,��3�6��gV��}Vm$�v���u��U�V�x8��v��ܽ��?x�|��_e�)ef���`�	֒�S)����՛��ye� 3��v�F����W�Z�C[@O�ݟ��
K�����HTT����
?�iR������`�#�a��ӧNs4���2 ��nVr��ƥ�Y�����iz��[�8�R�j�2����j�z'�����0�ƱM��
C?<�l��qɋ��Bù퀇��ꀠP�P�)��0Rn&��������Pm���2f}G{�c�l㶁�2°�Sn ?�C���)��mDg'@N˦�N�Rf+ 9��a;�q�ח��o��'��;^[.�N8,Va����������s�4$vE��ٽЦ;jU�a�ߖ�ν2[����{�.'�ϔg8Jo`H��tу��1��g�N��^�~�dy��}x[�4�9��<J���H.%t��*�)ù�����ک_1A~��M�l`{�uD9&;�~���7i �?�[Ъn��r��Un��:���9��g���/J3H,�m��nJ��nֺIx?d5�z���qi�
Mf��B�1�;�0_�J�`��4=x���SsP�Sl��ʇ��tD�ä�]�_�kx��t���O��j:q�wC�@����A�m���cA*$�H��Q�?�H
���/�Vx����Ӻ�I�L\5	ްc��P��B-�V�:RH�f+WH8���;7�]�B���6����t{6k��躴�Ӝy'n�
vo"marZ�%ۋ���:���}���o��j]|A�I<��h�zb���ڵ�*d��tP�]r��
�
���#|`%t8ƉkW����/|���t��=�˞��N@�p��w7kp��/�Z������Y����x�gq�H!�HZ��p����������o��/�S�cs7 �	3�H����H����b'�D�mh�<��]j޿�ޱ3�뼄^G:^�P���z�*'gKl�BW�k����4���^��Wa�f��z���<�+��0N�����\�0�p�LJ}0���>�*$*����̈s��A��~�GQ@���W�ണ�3��)E�ж0��AZDpR��3�v���,V-�A�|
m�=k�K
�6�f;A�L�u]V�����洝�Z�!?pi@�^�pp:���I����&,�]
H�S��=q.�Oc#AP�����G�g��5��=�׭���]>��.�/�V~�3�0���(�<XpF���h�@�౩�4t�'V�8����G&���]E� �I��&	�j�Y ���{���w�vFE@�v��*�{w���\�[���P���ӯ�Q*�0X�+�߷ӭs�����O�p�7L��4W&�fh`��=e`�s4���
���=�<�F�F^��,Ap1Jj7 Q�����uwM"*����ү,ѱ������W��e�(����-�Iz5�nׁ��j�e_7�Q8J;��Ֆ��Y���Z_S�[!�[bW�7������@+|nۡ���Q����v �]����%�X���U:���J��i�I�A�*�ƾ	N6y�U�
2�7KT"��#���@�P��]��IhVVfx���]�n�����G]�wN+W�����}����cA�|����ɛL�9�w���Ĭԝv�%2 �CG	��J��L%�D�����=<�c�qe�0�tH̻&%.�HD�f�Ž��D��S���z#��j�ג�l�c��2꿴�Ƭ�Q�������,��W؉;�e�:�W����ъ����i�I�r��%� ��桏��H��4
��� qO�����uJܼ�Vn?ݿ�q�����S8^;�(��ߖ���kQ��;���YL�Q���j+i���MAa�&��$�Z7�x�E=s�n���]:>�eNხy{�� ���~�Q ��t��_L�T��)�VGz�H�=���d[�����jx�~�/����5�S�zR����k��Ҳ�o�:��nяЉ�G� {�қ���[lh�73��B�Fb(��ulP�;��+�bw��ַ~�<��#�{��/��D2 #�p7��`k�0ꥪ���@��-����p^��N�l��3�I�Y��=�˴#���*��P~o�J%�СY��e�YbIj{'�����k���)ѻbju?B����_"��!A���V��`�kѵ��I�Ԝ�(X�_�t!X^�G+ѯ��߭��+ׂ��ח�	ёSL�5��'�_/O?�B��W~AN_r��0v �
Yٰ�Q/��o�q�r N�����%��:;8!�U4DF�΋QI2�V,A3�U!2��tHa�򼃁�Z�sPՌo��CT�����������{
��*x�!��cU<iG�+��`5�����F��ѳ`,]�!wOOo�� Y�Чۃ�D?M�N�g�6�(�:UcBP����0'K�hF��VGY�����v����Օ2aP���n���7��1�3]i١Q`0Uj]jK����^�@AC��}b����r���E�6�J�GS���2W�+�a���i+�WZ�-��W���uK���Y��]� }�"ǹ�L�z>N�/[��n@�0/fo�b�K:E-w�����W�Y*s�)�R�qb�BK��<�V�[}V�x��(�$h۫Ph;7a{�vT�71�)L�2;�?��\�	F��>��'�$���'l݂`�m7�5���n��".���9�ZA��b��x!�\U�����Z]�hc\�%v���I�\�F��t8�S�+��>� �P�D�1= "(�z�r#t�]�j� ��R.U��w8֖��[���WYdt]�����=�~��a��ksda2��0siD\���b��z�_vm�l�oe�f��~�(����Ȫ�ڭ�4�V� i��[���رB�0Z�ⷈ��վA��b���k�D3+L�{z�٩߻ᣎ����B�;���ϙ��U�W_w
#���-��kl�w�.�˷�5=��k��X6n�4�5�럿4��ʀ��q$휙b{w�y(1,���(��V�k'ϕ�0�g&O,��tN�-� +Q�j�������OZ�%��[������ͽ��6���������m�Z�6��n��A�X`���s�i�3,�m��=�J����Yզ?%F�Nk�m��쥲��4fo\�0�D%w���&19����&�:,;$i�PF�0U����(�ei謚�+j��Z��HPI���&�b���ϪmvƉp��LB�K	�����5�*L����s��f5em}����˶�ce��ʎ�G�*�b)���5�V�-d�{P�g���bd�C�j{,�$ϧo��2_�\z�ϝ*���$fi��[e�m{�8��r�4����`Ί�I[�>�]���2:��m�8�uŬ��]�o�(DP'\#�-T����b�����20#d@�3<0c��]Hɴd!eW�ˏ~�ly��قp�	a�K���Q@b��V	M���_.�<z�0t�%�Kp�A2��7�����a�&i��_�����ұ�̈�s"���=��@U_ECرc�U���<��F���M�҅�e�v�I��N��
n�����<�d�Cv&���_�qy/g�G�;��B||:�PE����j�2�@ V� D��AW�A�'́�mdH�E8�����'�Q[PF��-����|&QWK;m��c,�`���� 2����_-��O2>6��_�>�d����4�r߸�=�I뀷�4"s}ī�[����E��ZisIv^��eh�؉�Э�e���쩧�5��8�{"���)h���i�K�S�!��N	����?���S2U�6��dm�_	�W�$R�����"���m\���-���/x��W
q\s�0��?���J���W�g>���=(������k�s&�O�U긦k�)�}�N✝r����W*��vvvjYuݞ{61
�@�%����#�s|���"����!0�RpH�FX��ﵭ_{��<�j�4.9�YW���n��~�]������TG�-�p1gf�����C��>��2�O .r`�m���fv�0�90yj%���6F��^(�{�P�L�2���rP�1Jl	r��4c?F�M0^�7��KFV($�p�5F��Y:�cf�#3.3�H� ��9�,	ڼ���M�@7�[7mSks(��Q���fZ�Q�ݱ�ʀ��:��hy�C_,{�;�}��&C�#"����Α e�b�vR>�1��X���A�Ñ�,���!0�{ �!\�������se��r��'�^\/�v?R�����������X<z���d�A�2�6���\B��8��wi{�M�C�*��ܡsq����D`���D(��b�3��G'C�>��nK��L��8��GF��%k��: �9,��������B���]{=b���K$	D�JX��{�����./͚0��pDuU���0�`U�x���$E?���O��!�"�..�2ki�-"sWf�F9:�&ߛ�k)2���s��r�#ͮ\Y&��K̬>�^�g�:�z5_����W��%�
�P;&��k��3T,27�b�uz��JO�!OAꒂ¾2(�G� �Dݙ�(ɧ�ò���%�0�SG�����:��Z�j`� ���E¦D��J7�Π��60��1�@����3���nw_\+���K�~��p`���X<�n�0��F헀;��F�a���'sJ�aZ��~��`�2L)N�~�`̜G�}cr�}eh��Ց����ëo�}'�+;�͔�;0�c�Qץ=+6���S�:εi��b]`$5�#8��I���o�Z?|�M���OBދ�-
���
���֠�貴�J�gX�܆�i�:�%V)���/�C)����~9yF�1�LL'�����9�ld��q$�{ \�܆��2Vm�ϰ�!W@\���@��0p����O"�?���I�*Լ�5�[G���������L���[��K�o��L9zߑ�q��1H��U����$�/>����(g8#4�;� � ����u#C�9�"44¹D[�T����3#�PtK�5:s��8�0��UņZ��E��rq��.C.s�sTg�� ���A#�@�T(�8J]	%��$t�|��[�n�g��6T�!4�����P�.>�T;���}G����0�9�~�;�)k��x��ŀ�Y0�ɰ�/-���;r�B��Pf������0�zlm?>9P��88�W>��~�\>�\��|⻮ܓ�3�}s�e�q��m2�F�סLԕO	{�)�=R�������!�6�;�e�,B�;M�G�]a,���&�1	�+���=<�R���5t腋���WO�*�'��?:]�N�9�l��R��@,�p�t�v�&�'����z~���%H2Wz9��]jN�g�� &ma���/�G��	�������:�����*( zp#ҙ3g�x�U�m��;y������ˣ�4���d ��3{اq���?���	հ���6��v��2w�`��*l���!���v�R���Y:Kn@��=uk|���\�T8�荩�`�j*i�՝;��ЍJ��&B���Z�r�aEb��Ce�՚y��<7�M6�]�Tz����>�}b�v�@8ćN<�����nd����2�R�0h%2�@�4���7�F���>�����} �3Rμ�b�z�uV���2��<�����G?��������<_>����	�n���FI��K�Y���0��{hL��LԞ{|@0�F�i�Pf�T_ӝ��g�j�Ϯt�\��i�&�FC��ی䅶8ǊK�,k0y[Z�
AX�X��\���s�)4j��|�5�-����	��	S����\�<~$�0��~��2�GQwE���%��lr���[�����_�g��}6���٩o&�@�Y��n�k�k���K�.���$�I:ш�vRr�6��!����Vi+|ľ�%��S�����ag�Mu�h��{f�s��33�Q��!4��v�F	����3��em]5-��sU��"h\��:�uE9D���2�D�פJ!p�G�F#�k ;U4n; n�c��睚:A�J�ʒqhϥB�=���ϖ�*?��3D�~�m�ga�[�GN��)�BV�c��`g�*}��:���p�ie<�N��P�aޕ��B0�w*?ҭ�O�j��\��m7�+S㏖�Cϕ�o��˫/<S~�7�(O}��cO}�<��/�2����q9��~V;n�q�� �!VS������l��SQx"��E|Y�5������پ��	cF (|�Y2��f�ҩ·?is�A��cSs~���a�q�JzC���q�v�>6v�<S�w� ��x��T痪�B�:z�Ƶ9�!Ű�"�/���r�����l�4�X��X��/�hd?���|���Dp?�m9��@�;����lf��l3���;SC}~�`G�k��i��g��	
���1*�]�Z�ݷ=����j�g/��5�۰\���<��j3PX����� 87�pU�"DTEō�B%�"d�B0A�]m�
�"iSV��wMN$(� �7�R1G�2���U�����Ǐs���2w�5lL�Gl���];�T�VVL�06�T��y]�ٱ�-�p��bXf9����p63��/m�iO�^�����	�����1~�q�LZ�����l�:�Eq����������7�����㏗�����|���iy�'�i�5�t�}aƕ���W�s�iRB/ ޔ"��/���*����}���X��j�1�ډ�ºs~�7녃Y��T��n�~c@1���Ǟ��� �::M��c������_������o�~����ķ��1��n����W�4Т��01T��Q©�S�u�L�?�?}L�m��G[UhF����)u?~%���o%Z�&$���g�� �i<���"j�^���D��GYn��Ɲ�n���Ӌ��vs��0��S�8\������D�@A@���a��5����!*I!͸F��RPyPٍ���c(�ЄX.3lR@��z�O!���/#Tn[�ڮ�K��˧ʃ�<Z~������o�g����t?|��ݺHKL%.�1�#|�����r��� ���2�U�?��S,��BӺ̖b�`�݁f����QƮ����74v�'.��15s�l��0L��LaӸ�hT�1�-��,/=�������oΰR4P��ȓ���ʳ�|��<}6���ߗse�!�>�1��%Ia��"r��l����n�U+�`�
q�EO��9h�����g�V�3c8K��|�ÞdjV�,�J����={w���:�`_���w���@�@H�U�QɶO3_�NA����U&X̉�O �,�\����F�P�w��38�;����&1�+}˪���O����<e������_;�\9�F.�6S��ГS
|0 ��N�R��� _��`��Ò���
Vi���"�]I�!4[��[? �8;���%U"�B�~:L����>��Qka 4U���&=��64x����g�M<��_}����8��0S�%��q��p�~Y�{߇��)�Vy�o��g�-o��Aٵ���ڈ���0��"��k�
����'ڏ48����NVD8��e<������e���,�Wvm�]^���&�h���G3Y*O~�)�R������w������3���'�K����W�����嗉z�<�KOE퟽v��v��쐿����
	�]e��w�&�����Ea��x]�#���v9��0�3X�B�Q�>^%����l����
j�X��wN�ӷ��2�5v�
)V���}���W���ˏ�~�|�Q�� �M��I	��[�����xXz��
YJ�j�;%(%Kl}����V� ���o�|Cu����N���m���;}
Kj{�l]���o�[�����۽'�����?���������>�{�h�+S#@Q)o�`?̻k�4*��m�V$2�۝U5+��N`Tu���S��q��!��gY��@����%h&��0BH1Hv��%�u�q' Pڣz��e�s<���ū����~��������>�-�L��ĺ؋�a�&�,1��r����ԓ�.�<��a_�y�2F�%V4v����'R;ܱ1�C #�S�%��]���{�Gx�<N�� ��r�]�/L���izp��\~�\>9W6�A��Hy���7��u�ļ�YVF���wʍ3������?���S���~�|�/���r���e7+,��Ωh��9�Y9)ZV�����8�C�������;i�
fI�d�W[����7��w[��a�p��r��u�\�c0(�0WC�(xލ��Ј��2��"k�Ç�g~��\�p����k �?��_�0�6��M��dy�(�
��'l�.#+�&�m�d�7�����^�\�|�I4������ᡇ�c�q���p������&����ɸ^
�6o��YA �kw��w��&�Uo�'��nWkq�kj\>������!bkZ�ߥW.,�)��������>�4��r�@ʿ�}�P�ԃ���gh���)v(��gϼ\~�����/�=��s�؁�r⁉2����D4Ze*6!��i�%(�p	�e����C|���L�&HYZƠ���9��n����ʑC��4(�z�|�u��������h�j����?��z�|�׾R�����?��f	�3���FCW��w
/Pw�kg�j���
�6���.�����V��;ue�%�!���
tz��@�����ϳ�t�<���o�#Ǝ2=yir��\�6v��3��K��� g�|��8fU=H�Q�J��o������|�FS��m��fPմZX1���@�uWm�^������{s?!9���f-���
����}�w�S'O���je4T���X4z�'�ϲ<���3B�@#N��T��J��R�� G����9( <���Sп]�Bb�[�^��ΪHg�F�Z�:���%NHD��
xϾ���P��/}���e���'>����g����K3*�N�	#�z�ٳ/#��[V����#�ʱ={���β�ֵ�R&�JQ��I���	�.yz�\����H���Rtl}{�U�܏�~�2�{gY��z������r�Ў29�赫啗�)�8�}��_������PΞ}�|�O�3�/��}�%�I�v���OwK�xK
� ��/��f���.X���s��"�w]���C�����
Nrx�2�{y���qkG�?��?//�	����'?
PC��� ��rFm�]����|�i�s vK9�8��ъҠ���R*��>���x�Ž�x��X�a�����v��L����N��0ˈM8�qM��f/ޕ�d�hΨ�ի�&��V˹s1�����p��K�!`X��yD�	l�8� �4�<j�Mi5<����E-Ah�iId5-W���^�U��
���PO�����ly�*�=�x��w�����ޣe�y�Bj�<wo+�vm�b�)���9�����hh��)��M�Q�C��V �~N���)�cmĖ�_�O��.�.  =Gftb3 K�0�[��/>��:�&�'���^/��W�\�Y9�*�7��O�A����-/�x�Y�&����Q-�Mn�1#�4��>U�u���m�Dq��>ו�>�		��w��>���$��j��!� ��c.1���B���[�~�7��<^���o�^����K,��� ���[elj���N�$r�Q��m��8]iG�`ΚGYw>Z	���""�X~�!ݪ'�t�9T�ۼD�x���;Q�WG�}�S� )�|����0:�� �E~�{�zs������;�R���%��w�ݶ}������G��?.�A��#�V�%�Y���WX~���/و�
!#���ҋ��=���7��1�޵+����1@���Qߺb�ᷚ�S�0D���	Oͱ�a<g��/��'��t۶M��Mc�M�q|��jQ�t�ؿ�l��^�t����)��I9h�6!������g~�em|�9r�U�!��?@ ^(�������+��ʙ���L�ɨ�?�B 	: Z!���������:�f%^V��h\c�������`�CCn��s�x(�.������K�f�]Y�_+��+��1 ���f��P����y�-�(`�=�!��W]�n^=�V��M���g�q'.fc_��W��Қ�	���+��ޏ u�e�1���j�j\�^	2����?�c����Pš
�.#�gv�DR�¹��{;S�� Ƶr�ȑ�|�0�o��z�!�4F@��J|[���~��&�2A���x�MN�k�4���\߽	����0�L����#U��3��.��N�p�š9ڜL�Ӟ�s��Z5�8�&��ڃ��:��p��~�Ѥ F�� �8T��e�o�:E�WC��%Ҷ�B�P�;�ت�da�3`��c�Ϩ�~���̊�N���_-�}��Q�_����f�1�L�]�W����w����\;�z��f�P�_�W<�}�0f�w;a�q3z;NO�,3�c<>vt[�VΟy�������ʯ~�|�7�R^}���o�ϛ�>��-�����"Z �!��.Qo`_��Y��3�荴M���>Q��?���)�m�{up�x��:��}�K�)T�_�C���Fԯ5�R��*���W1��Ĳj!8Kl�<FM�����s�|�,w^�|��I���J���-�����!��޽��l
40��26i�~S���v�:��Bｷ�K��}n}��������]��0t/�sPs��6�'
@B�O�Ĩ��C�dS�!�0&2�ϢU,���2�:[�%�L(Dnӗj��E�'58�ڀ���Л:z9b9��w��F��`�>�V�����J�Z�F\���NgZ�[�+��i�3��>p��[����q �����	�c*{�)�Q�W0:bGܵwѼ���m�{�j��
���|���h��A���%C�2��x�m��*���.t��r�~5�������΃���)g_�Y��W?�G�����lY��� �v}]���2��W�:�
��𨶇�4,Fc�k[B��{K����}.R�!1,�>�S�J
,�8=��2�G�Yw\�+��� ;�2e'��F,�-0݈W�P'_;�>g8��������M-ښ������c�l��������ٽ�y��Q4F�E� z �
���1����lv�ʕ����`����U��m�y�Z�-���y8�q\��\���\ 2*2��3R�������^jLg}��[�dM�ڰ"��OO�P�j�"�R���O���+�|�Yp��E���2��Y,̢=͗��N��8WN��by��ɏ��绎��u����_���޹��b@Ʀ��9�0��W&1�>���ip��?��?�����?X��,��W����o�vYBP\<�\�|���m�jו��e.�'�L�*O����l��77��Rt�Q�t�ihu���Z4Eh��gޮj$�^�|�����X�uRq���9Ծ���&	�]���ˋ���v�L�U���F	�2il��>i���lw\" е�V ���r�v����o~����٦i�L�w��$b��|'#�����g[.%��4�Vn����k���ԇ�险�"$�P�p�su��2��\�y�0�n�ҥ������j�Fn��6��3Q���}�K�n��1����E�l���0��f���by�tuU<�5�?˓��Z,�嫳ؿ>Tn��c�]�{=)la�C�K���Ջ�^`�m��U���i��j4L�=�B���*�*C	oKy��ѝy�w��/L�Ng"�Uq.��e�ۦ��H:�R���h9~�0�)��?)���-����%�4��}��7��{�{�N�:ò�M��j�/&��]4�����Up�'�%~Ɏޘ�$6� p�/���)Z92��+<
tSVJ�+�S6w�1]�y��RN�8��av�%3Đ������t�/6!#�Y�-�@�(�h�hm�|utrLG(vFK[C�����=F���~����g�S"y��=��Q$��*d�|��X���%�Ndi���/�+';^��v�#��ͳ^O����������WF8 @�ʎL�(�Nԡ�g���A{|��9hG����͵.7��%K����-沍��?lM���;!�.�'����Ѓ��}\8O�&�x��a�K�>�A�r|&�<6�P��Sa/�ڬ�����nS��(l�>�@�іªF���Q��8�i-� 9��hw{��9�}��_�z���h6
<Eʿ���#Zݱc�ʹ��ȵ�f��6��HZ5�ڞ�aH
����G5�V�@a.������/J�ѱ;e��
y:M������ 8�,3O�4��c@������:��ب��n��V8�o�݅�Y�)��u�A�����������1gT�>Fm�[�}���HS���^��.����ZA��>�>��b�a�i#Z�%x���\R`o���hw�U\%0���N��㔤�� ��(di�#���v�u߽~��N���+	Häe�X�@)�ћ%Ԏ&�x�"u�	�=dT�ld�  @ IDATh��'���	�J��!��Ξ/'�?Z�o\ŗ�S/�[7�r��,�Bsx�b7��
�+#��(����N��<�Z�����N;��)��W�����SO4-�u�O���Z��ڛU0�_d���>W>�؃���hۿ����|�7>[8���f3ӿ��U>��'0,��+�/�y��3�Z����~o+M�¸MB�n�u�
s�Z�E��&�����gVK��x�g'��K�_e^lϨw��z��KC۸���o���r�$����a�(wj�!a,�`1�|�e]W�0��|���2�s���6ד[��"���hj����ڰ�f}����#����$�:R�>�2*!;�9�eG��|���""�<�V����5E�eP��UC.����0s���@Q��݈�Z`l��Q4K�e䢬04�R�NH�	w���5A���q01pk�Fy�����r{�$�k�s>�����7������k��,GS�t��S[�ڎ۹�Y=<e]��?D��=m�wb0�yՎ�_+�]MȦ⸪��<m�m�H����u
Ap���Gs�%Sr����?�J�Φ�_|�<���[te�zY 0�x����כ�PW�����T5��?���L?�Mu���`P�~�C�yШe�ڃ����}� 21^��x��@��(^{��v����^�g�U�����_���f�Պ�)�U�0�IP6-k�~�jM�ܖ���a�r��6�5?٨��߼�je��T+�O/��Z�,�[5�d�Eek��2m����~ӑv��jj�������!�6hԳ���� p��N�T�,.�a\q`���0�r�
Z�x���P/n�\7��8���8����ዴ��%d�;p5<���T�� ���B����$T��_���Z��T<�>'��K�������1ݽI�7�{�^>��O���@g_=��#1/�_PX�b����wϔ�{XU�͟i�����y.�����ԍ�&���U�Sc��I��\��%�u��}1��� ˚��ȩ�#�s|i�hUD��HA������q�%d��GP��Q��G\����c_��/.S������x<^=�f��M|CX��V��v�J��*p�&�i�I�8�ى��\�W#��\�)+�P�S
ϵQ����1G�IxI�q�]e���D�����A��8�If�)�X�]�p)'s2��Cn�/�r
�ޑ�u�Q3a]i�s
}����kX��M��ۥ�Ʋ���~.3'Uf����ݓ���(�+D�7��L�F����bx�HPzB�������I~��D�r�|h�M�D�����B��pa���`�5�D]���Xv·B?�a���&.��2=��Qv_0�X�EoԞAsS۵_82�=��^Fح"��U��gTn^�T.�;[�x�d���e�$AiQo��R�����N��pi5�&�$�U&>�ZO��R��m%G�A��*���v�Q|5�)x=�Ѐ�uɑ�f��l��A��q�������hl��/��������"�c�x��<�\8O�Q�R�/ê�+C�(��Ѣ��ó�LqBk��֍�i��C���6���yՖ#SR�
<ʊ�U�rI J]�W._d4�Knb�N1.�]��F=�q�4�2>0���̴�gR5sI�"�΃ ����w�����he��r�G{�}�@%m�O_l���>����o����{�k�v�������
�ӊ��X�oBےD��7AI�mY�b�a\s�� %p����ڍ�ۨb���\���B��Ly���p�*=eJD�G��hE��*�ڴN�>����LA��\)v�A4+������!Tt��j��+Z�.�@E�)�^ �o����F�0�Zڽ�w�y��՘R���0�p����Ap��JK�IX� �e�:���U��I.�2��gW��h���{�v����Z�Q����ʸ����g�i�|����m��[� ��Ȼn�D{qJX]�A�B`$Y6!��*�J�]�]��>�s�]>Ս����:I9��/�Xw�n���Z"�5�O�z�R.�8�4�*ͯ�?v|�1�i��K]��]����Q�$���7��Dp�����@�Q�����lw���hl�q��њF�#p��H������|�:�g|��B̅X�Gbi!��5:o_a�hO�\��b����W_}�<N)G�޻��)��v�g/FV� ���� v�?�]��o��8����45�_���aR�����F�ѕ
�ܔ�����2|_�9UhLgw��F��;a>3c ^G;*	\V0�a3qd]~u�zࡇ����o�8��,�G�LON�Ɔ�ٛD����^�1��1t�U ܝ���v5[�}����/G��{9�Y��x�ʌJ\��]�x�Dٹ�{��t����r%�*�����H4�����.��̻n!!iY:O!�ă����ĭB*���_Z��nCSś*�O�6��>�����A�ݿ�M���,�"hv�ھ7wX��	a�l��>{p��|uDw�nr:�������U��ȶWBFq�#�k���}j'��Dik�B�J�z>갤����!�5B��l#���;���L(c�t��H����T�l4vV���u
�Z�'c�C@�'d	m����w�#5'��b3���n߽��Q&s��e���qs������QA*�:A�O��a����ʵ��$�J �v��#����C A�ĈXgd��}���9D+��Ь�#�E��a�=��i�e6��e�c��%��v�\Da;�ͫ�t�Hۤ�"U���*p[���A������9鹻�J�T�o����oC���J��h	8۸�n�i#������cŶ1��O�_�P.��6��V�v��K]������;k��EJm:a���Ĭ[�������Q�m�ݻ�q���0��H�2�sy�C��S�m���m��(�<�/^�~]���c�S��=�
�8q���� �|���w�9.�;��lW#9����"�i���:�/����s���3���j�q,f�oPc� �y�m(+�S�����5�9��_���_(��]Ld��m�a$��
���4���ǟ���O�IR�Tc /)hBЅ���'B��A��Q�=*9��د��h/S�q�O|��G4�Q�@�-:LT�iڪ�V��vj�v���w���Z/�?�"W����U���*�Һ�F�Q&�3���jݴ��:�栚9�s&#����3t�R��f���DAAj���~ht
k�#��;8(y��8p#� G��%Y��0���Ӧ�����פn�� d-�e����zb=�V{�k7�~�$�B�#�Llr�v� .���t���$�l�׍�|���g��Dc�C�Y�KC�gB0t߇u�n�%�;p"\=�����S��j��L�hش��UU���p:���EէC�A{`bO�א�~DT"V`��g�M�,M�ľȗ/�}�}���=`0�c�Q&J<�t���.:��3M����h�(���Fe&r@��,��э^еt핕���2S���������F0U/���/�X<�=�=<<D\C�0i�\� ���!��$Ѐ���"�
`Ĥ���h�R�.�q�q���~�i8B2H%��
][I��IB+�	J�'"�0��"a�vx��ϩgƱx��㲽t:��k� ��m/���I�K����{!emFX��vF�	��w�~�/w�����!˯e��œ��� �7���{D��ƈ%�^�D�`=�X
%�T8��H���go�ȯaCQz_tw�����1�w.�i�\�2��W/Pld������䬝�_�B���	��ˤ�6�;�Y ,�]ncbafQ?�Cg�f��DL�oa�sg��C����vX��Q���tfs_��D��I80Wp_}�2�����!@�0��5�R"S4��8����s������[��en��΢FP�^��0�a� �P��l�3���'8%V�01v4Ҿ���~��orL"ۮ��$~Ӎ_����2^��6���ˬ���	�I'a��Ye8���Ԁ�4c�{���Q��
nP��>�����*o}�w�W��~'+n��tR�I�;v)�|�,.��edR>g�x��iE5�ⅇ�^��c�5��L� �McԺ�2�����]�w�{}��Zצ=�lf��,#بs�3 ���A��aa|���֙N&A�X��:����R�N���vV�\��O���z���3�>���RDj7q�L~�@�#lL!9� ��:���=K�{�l}��$'�)������~�5_D���l��ђY��X��0�*��gzb��m���G�T���KN�1�xE�t�5�s�%*g�,�>8�펅�I��#?B��)�6�9��JG��M-���$�S0�jp%$)M�ԁ����ܪJC����ρ�y���G�1q}_b�����;�B=�����C���<���	���x�����L�˰Yж�>���hm�I;Y	x8�o�?�G<�l?���ɩ�+�i��Q�r ���f�M�6P�l�%��΢*^x�*!�b�@��EWi�+�)��Jw��0:�z���ƴ-�I��O��3|������/U>��+�@��=}ʘ�Z]��89�	[�Kg�������@αqT�Y�ޔ3t2W0���"�����^�]0�J.%����@��������̙:���.`���K\(�ࣰit1���1�s���+Uc`��X@9�d��|&> ��#��,� �q��;���'s�dvѵ!Ϭ�A/g>�[X:#�F!��nS#"�!W=��� �ٷ�{���o��]���8V2�����{ oP}(dZ���d�����F�^��)#�%^����s���:�<����i�PŰ�2������T������N���ݱ��Ol{7���-�,�u����Ƹ�
���d�e���o��ƭ[8I�7�\��A2����d����2���-�����M	��d)�1dw/��CR�Y�^ ���;������J,/ab���ӝ��D�C�b���)�')�-�<�-,����`,�����g��.x6�/���)&>Og��)Rw���%��̥Z%$g�J,�����l2�:�ܑ��is.~Ni�s���#)������Ƞ�逶��a���uvgO�I�#AX�:�RKx���6Ć.�	�v�������ڄmtGox��z����ė�|��bvQr���5gZ�X�{v����s1����NbHX�(���4���$�����9ð�K��s�����+�?ԡک�����^�F�3?��!@C����2t�C���^�Xq2���LlWx j�[%�GHU2#^h(������`��;?��Z�'OM�O���G�'vr"�/q�x�	n�����*�}�K�ʕK����a`E�6ey �̣��ǐrZ�eW�L�W	T��S�3�z�H���HӾ�Tѵ6���V�vL�:`/Zn%�n B��T?��Hw~����AA�6aw$�������m��sR�J
c":�&[�3	�'g@�D����Y�%'9%�X��R��.�!�'0IB���̪D�Hˬ��TO	���{��a ��Q@������mdi���%\�RN��pO� �D�V��8J�}���Q�<��I�ۗ��K�C�M�}B���HN������=����h�c$��8�|�#,�u�d����3�6��_�j�FV���?�����c)j5��?�r�`/�2�fSm�x*"A�a�P��ϲ�*0W��lK����SA�f�nDDc��%M%�	v���a���ʵ+�� �)��p���믾/cQ,�W��DY,��}W9��&�C�G����O�:�%���a,�K�]������T�\���<�:�E�y0��(��98L�u&���}˵�0R����~�C����F����2q1a2�ĸg����� ��q��jf*��[!��!AWF�hפ�� �=̊��9�?�F|h���K��#�@TW�5���T�Ĝ"�"b*ut�ݎ8��Z��bC�.g���$�/�C��Wü'sS�P�|9�u�T�߾��]:����l'�F{LǴ9�~^t"��j��-<I9y_�f>�W<)(uݥX�D�r�����ؕ�����B�bj���.�E�̱���8�(Yǆ�T��9VҚ��^~pD��ۍ�i39i��3�U������)O�<��Ǌ%F�\]+�ǩ�zq��Geb�hE��"�|�""�8N+˫K��i�.�g��X"*���M�F���V]=6�,�����N�t��Š�(L�P�`�|�^$���@!=y�����}3����LC������-�x"+sR4�WE'7w�����$��v'�u�8��  �(9H�RS9uPt2?%ʓQIZ�A%~��B��M��Cg6�9�C�3&,d�t$���*�QO:8��I�a���K�Vκ�j��?��^�'��AܬbF�������"��(�q�0��ڳߖaJ��o�A��gJc쨯�LTX�T����Fe����d�L��ҧL,W���,˞���h�l�03F2	�0�����w�Ʋ.�b۠����G�����?��<6��'Ǎ�),4e��C�: �`�h�HD+��9*�ϟ�)�7�xFG�d����`FƦ@�1��f����N��ɍ�Og��UD��%�J~��$��y&18@4nW ?��KސT��*FwQJ��i�m�~�}m9U�&Y|��X�-�{"m|s���C�;����f��&m��t[����k�G"�
W"�C��p�K�f�M��+ҥO��w�y�|`�9�R�>���Dh��**2�^0u�'��-SBz�^φ���-�-�{a� s��]�~�$ ?���~�7C�c ��}�Ǥ������/�,�ZwW��ײ$d��e�LJ0,�_B�K���O�A�iH?�ߴ)�����?�55+�+U2%�Ah���e��^n�s�BJ��'l�J-ۑ�}��ҍy+��ם��}���N)��ۆ�tM��&�^T�����}7�l�\�{(@ Z#R��,����Ys�4m� j��'.�^�R���n��^G������|��ħ��/Y��h�%�秊�������tx�usp��,����D�������9$�?>�;3�!�=��2�Jˊ"�"��%�wc5�"O�;˪�c��.���Ňkg�t��@�H\�!�9k�R��~�4B\�W���Q�����ŷ�ѴC�n�2�J�t�-,הp$�;hSL6�xk�����z9��~~�1Pv��c�D��  ��E�Դ?�]ڑ�m��l[����>�� ���'W��Q�a#���~��������&�E���6"����<��虒	�e�q$,l�;�C5��!�����XRQ�[X� ��"[��"_{�5�v��pm����K`����3e�8x��/:}�݃�D���m��Srt�&��c^g�ܒ1����� ������1b���Н����F��Z��e�~L��*�i)����D�v�GY2����1�0(��B$Dz������f?�\�y�b�ԠO�,{<������3���μ�c�:c�b�����hC�=�-�	#@mt�c���  ��A'\��@j���A�K&��@�1�i�]Ѻ{L+2�"��;H�>�Ĺѯ&9gs�~���P&��pB� }u9V�
�X>�y1�G�����-��uX�7|ȯ�q+�^����_ǝ�X�<���<" ��T2J?�8c��i/6Ȕ(�G&��< ���K�)^0�Cb]l�ߨ�s�=_cgw�qi��{��k|,�r��N Zl?C��v
��Ʌ�:�?� � |n�y��.����i��J�a@�jrVP����1bh�p��dTk��<���R��>ץWD�2+Sj�3:k�_�;L �S���L,><>q׷��w�<"�$�߁j�M��qȅ�����3�]5H�L<E�O���H��x�*�㒾��b�piMdP�ɍɠ�0��B}�`B3�+u���)�ؒYh#aFj3L���g¡�����k��ӖȚ6�«�i� �dx�rl����r�Z�N����T�/n���d���$.��i�K�K�ʾe-�BR�B%�*�xh�)���K�^�����5p��e%=�81OϜ�y֟��X�%J(��p�	XO�$*��G�B�Eї���>�^��º�`$�=۟��,a��59PK�A��l���ַ�V��>�pL8hXL���-�'��!dS�M8���� .�pBV��e[���1��R����@ԂPvPD1�]9k�_�7m�$�E����ς���hs��5s��Q6�y��bnf�����z�3��LF=���#�{̜.�ˁ2=�y{�]�̒�9��!g����8����ٶ�P1x�΄0�#�Q�Fu`������n�p%�{ϸ���]�L�7�AG���M1���7��8��}��q3��A��(a	W��X���09�k;l���ԧ�K�|+�K��#�5�L���7|u�B �L�x��O�=�2v��#����K�j�~&�4�
#�14�#�Qv�͌+�~��ե9<�?�~w��Z�`���8�\�R/��KW*>M(=��$�/��4��{����fl'����0��6j�4z��LCՃ�Tc�+L"��?���ny���8�DN��723��,�C�b�KE:�8s%�Ӡ� /F�Mq��T�CH
m.��b���+yv���	����J���Ϙq<�q=������P�tQV�s+�!�$X}Ο���˾�~6G1���e�B��qU,N�����*1���]���O	���HK���O5�ՙ�������6/��xgt����{0	v\&��LO�M��)��׺��PA��i���!��k�����0Ex?©N<٦��{�P�Y�+,�����5O;�p� �4m��@��R����!��T�`x�K�ea�4�!���')����ݹ�v�	�b���Y���ih|�Q��˩�n:�c����J��m��Q����R@�A0E�B�?�������%�)Fbh<qPܲ��� �Lbzj�Y,�U��e=g�h	�8� {���6�RW1~O�*]|����ӕT���i�>�����V
��wb�i����{u���2�j;뷈��|�u���䎏׾����`�8���pN��ഭY��|Ʊpj&��]�����1���S�y+�y���c��S��@l�qEB)O�pe���HF��sp��#�9!^��P�����(�x���5�qJj{5�T�qT��p9^�H�C$���O�%7�bH4J>�C|�z�qZWOv2�2D�h���4
V{ږ߮4(��
���"����1����O���2mH/1�F]ݳC̈́�i%�g�M�z����̈���G㐸#�]���'ؒFYnD"����!-�w�V�H�=2��x�:wB ��D�a'��$��P��S�Sh���F���-��/�I���R "ś8�6�(�g�zW�9Uzjz
=�9�+ۍ0H����H�e�h��?dA��NxCR�菓1z��!�/J!��v����;3`�Yv�Ô˜����7��]g�!���K���	�ꘋ��q��#�)b;N�u|$\S0^�l�?>U4wYQ|0�Ӈ(��\�@�άT��;G����s��㫿�r�ĄFE��`��=�p�����3����� 2g�*	���#q���б�J�J->���M1<�C�޾��"VP�MeR!}�$�Y�O⅍��Ѯ����3�p�n�k�9D�`�J^ǈ�S�s�o�v)�.�otH�&� �8:2G�e���׮Bst�)�����1�(Qw��qI�^ze��|'�ȓ�br�R��/%��ò�L;V1��C��ܹWnܸ3�K/_��8��ɦ�A�Q��\�����,�R����pNK=F?E�8�RZ���=�MDOt�K�{�v��~����t�.��[,'�L�2�x�
��%�����k�)���9��L/��cH}��q�������b�2�p���f���!��|0wE�*�TFF/@����ڏ�w'�2�I�vׯ����ح+�#��&��N�-�^-�_~���qR���0����n��Fx6ބ�wԔuE�]���;ID�l�������d�M�B��Wp��"S*�!�V�>��~"/����]�J-�.���&�z��$�[�j����>#x�u�BE\��7��F9n�V�ZÎT&q�,�?�����c�X�fj�}q�W����6���0�r2��_�QI֕'�z&��ӆ�yL2"��U�TQ��b����c���r*�e� ���4ƽF��nA9Q�\�� /f\�a�����f��`u8��5�����Sdg��*\�7�>�����}��_8��I��"����ŨL�x�� �I�_�j��p��0|�R"���Z/�Hq�i�Nƴ��q����d��~0;�
o�>&'!u�.�]�t���8��-����m�:��� T[dn�|��f�C���#tv��UD�"_ef�I&����]ޏrrz���d��BB�J5M�DJ�b�}�"���,G�����[eqe�|�ۿ��s���D{�/��܍ Ól{��`�3�
K&`�`PO�j��s	�]�';��6 �������-�&�q���',���y}�~e�� ~�8���{?(��Yr!�z�����F5�;�Ԍm�o�rM�]��D3�p:I��&o��[���~��_{�:a�]o9�]�X��ˤ����.�S��Ia/���S��<�����)������kǻ��u@���O��$1;8<��
bG=�ǡv���,�n�ljv&A/�؏��ᝨ�� ��775��%%?f��]a��Zd��v�4�c����[�[�dV&���ոWV>�'$�ɓ	f#qf� rf���b�N��5N��[���;����F�@/'��W^Vٻ0~�u�&QP��Hʕ)Ѐ����@��������M�@7�o�l���8
G�jU/�sd�_��L��79�6��G���ynx�!˕�x�0<nol�G����^i�:�\9��p[�f�f���w�Ǉ����.�����u~J)m�H7\�u��/Q�M �J��c���^qK)�Κ�Ga��{�~"�ԇ��>��C�/��n2�T�;�n^�Q?$P��3��e�}�ΊW��H��j���KR�狼����׿U�pz��&G*G��X���z6��
|t&q|M��1�P�-��"ę3��{H5���$���@>��:]��Au؂ыr82A2�}��iI�T$��&��$��݊"b���v#�O�?B��5�1X+�mts���$�!��v� ��'�e�cg8��G�l�����M���L�~�6��i�њ6s����B�y��l���Sm32 	&J������Ԟ�b�8jD�w����Z����K��5�s����m���{��pʲ��+���W0�#��� K�Q���J�d
�vꮆ�l��_��I6]mk��'9�BH!�F\��㦴�uS����%r�w��1�N닫e1hc8�j���<��I�=��2�w�'��2XMd$��F�� $��nZ���?��S���}B�O�����Bz��ӯXG{V���q^c�#"C0:�y^��߂��B����߃����;;��!a� ���j����8V�Jg�A�@6���v�}��#��_��7=��3Z2�:c�/�&1�W� �� ?:1v5��*����o|�l߻W����<����箱�0\�ｇ��Z��ţW�����i�Md=�2��w�'_�}�#���A�""��jx�I�=���I4�By3��qs�T�Is)B����XІ�[�{\^�ޗ��­�m�Ys��Щ2<q�������+F℻&R����Wg��5k}�v�������a�:�I2:��7�H�b�:�/�:ڏ�I[���`��rf�n����Kpn�M��@U� �s�k�lE���e
��������������|U��� �2�^ ��5/=Zo<O�r7���\��٧���1�1u,]t�$jp0&��6�,:k0�!r�@���3��,�~,����*v�'����=W�^æ��B�/-g�6�Q�.���ˋc	��Q�M�!�\�DA�)�Rl�J|�{�!�hG�g%_�c��`����G]����S5�YJ��!<`i�J4��k��?
>( 3�#�q"�����[������Y�(Sl������',o�<=���kLA
����&�t{R找��bO��7��*'h��!:Ή���=�����?Ăm��A6�Qט�/��j���@���@�o�)vp�M]K��^=☻Ӓ��Ӂ]pf��4)�t��[�3n  ��ǽ��ċ���u�@ק��C�;�w]˩�����I�����O����E�'>`����C�X�a �l� � ��n��	B�+�¤���U�cʸ�m��.O{z�dD�D���i�N��
%l�g�X`<�U�v���7�m�YD�|{�G�]�L��,���m`m�v�&0��W������(qR	h��JG�Թr�����9j@�a	~�%@�W~3�:�Ҏ��H����%�`�_d�>8��NI_FqRxn���J��FǸ�|fY���Ğ�C�:i��9�C�{�o�~��r��Y� ��q�w/*���NY!�ܙ���������b���xƉ�']��v��a�T��U��'��F��I���~'M���C	��RE��,M&'GS@�ܡ�v}c�A+�z�xi�|��G�?��	�
���KJ`n��8��Ʃ�,��\��,��b���W'�i'��j�w�ꍯ�[`�$�ߚ�`^�	�%{?,��z���]�CS�S��e����y�Fy��k�R(:�"�&���/��	��H������Pzj�v�(��c�V�HF�6��B,��Ȅ�D
:���(h��u��w�}K����5�9F�G�3����f�7�/�c������8�F��Į�<0Y㧮�)��O"J��z0Ժ��k,��0��b�J�+��Ƞs��W��`?�횢}�<?��#�*���I�*M8ikei�1~E+�'��BuX䰠u�����Àz��壟�W�������?x��2}mI*�;���Ǻ�l���`�1as	8CcmfA�d��I|��g���8����F���9�r������$J��x�<��X>^*�e�<"�˙@�,��������a�{�.za�>=��x�ja	���Z}�&��f⢛I<�Yt
�/?�;�*�N@>?�O6�� ��Ǭ�	@��/��&�q��:!5�}$mH#Hn�"��҂NU:�y�j��x��d%CC�� tR���` +�Ԩ�SGP�as��HQ��@L*B!oහ��.�Ъ��_^\��[�HH[ey}���{xܶ�4�J�^��H8p
��7���2�iV���sx� G,��N��o���>�r�3
5�+3�$�{٣�B���1�r�,� F����y~)*���e��U��߆��hJ7����]����굗�F�ه�!mڈ����\���?�g'�o�L��ѐn³�qp6��ш��c���aï�g2.Z���r�Tz
S~ʠ�x��.�ԝ��:�����A�xQ������+���
.� �Q�2������]���"DEDEG�@|:UK����?�9tg���"hE�/Y�o��d�"�6,	ؙ���Ї8��n��(;8gu�F/�=��0>h��f%�DBc~��ƌ��@�!��(���"�3����x��w}�FJ�����\��܂����:zZ�D?���(*�`�=<z[X/3�!��I��K�}k}��CԬ�se�ԛ����9�$;̲�+,��K�J�)�[��@���ia(��T�$R��1o���+p�kq�� 
��l��=&ʭF�y�A�St�r�������+[H`}����������*�ҕ+�Q�0��(�:����=�}�a���R-L�$vi5�k�sl�B���Db�z҂̬�Y0]t[��ٱ +Z�A��Q�'{�|��7o���� �*���R�/|�L��0U6p�u��-���%47ڌ�0(��"Zx�#&:anqK��*@�;�d�62�u�s�
Q�A��kE+~�ky}�;nv��F�*q�2��!��^g��~e�O�Y�!^�}iDmw�|3�2�R^��GJ��P_��<ytO(�[yЃ��ar�-� ���k��c��p��f{��]>]�/�yD�Ph�z��f>Ĥ0�ȎTj���8,� �$J
gcЫ�<f?A)3a�bگ <��"�"��H���F�Ǝ��f'��s˭��,�}�4�.���Ge��9��	��2��I����o���Se��w����|z��A����h2�9z�SB�G
9���s��i?����|8@��[\�2����D�S��{(�˲���rX�b������xT�Y��ֲ�:�<n�;[=�������:�,��s�2pH��c�I �ʓ!��B��~x�GW��2x�Cm.J�>�l�Hc@���� � ������[����z�����-A����Ě\-7>���lZ)�O�\O�Ct�1JN�ΗeG��q�p�/���f����q�~��D���~�*+c�y;�\o���x�������+���̇kd)#�/d�A�d�4Jz�z�����eg��[��a��d2��A�8͛Y���p2���2 �)X��:�:�`2�df0�;�!ʦh+<N��:/8!��+�bQm��/̔����r����\�ʪ����ρ�c�{t��g�C�<�/���l�u����}������и0�҇^`�r�L��0�z@FDv>0�<G#�Vs��(�������Fd��1����֭H�*�˦N��쮓�7Y�=��`V���[|���w���������#T2P27`\Jd�̅Y���h�^>'rRmY~ko��?���+����o��'�n�2������ �8ˠ�b�)�/^Ÿ5Yv��<�k���9j�N95�P6آ��T�551U֎��Zt����s�P:�`@������6$-��?t�^�X�/.%�T��'H��/�|�������0���Yޅu���V������� �h���1�ad"rT1�V"(3�[��.��ɬ��j��
䆡L��O����J���r2)$�<b�ۯėc�����7Qԯb/�c�Qs��!4o�;���%��4` #8L��elDZr	�Rcsaɳo�kx�N�M��~P���C<E�p�> 7��ħW`6�!5��Ci@	�<<���.d�Di����3+�� ��I�G�Y����bs�A��g[��0�P�Z]||��4f|�c���g?.�,�~�Z9}�R�P�a0S� T�K�/ ���"�Y�r0l@�=W1�?"� �[?�%c�(hl�Oi� @��,IN\p���4I��H���VR<�8'P�Rc�6��ϰK�d�O72E\&}�uhQ� ��^E|�ѡ�э �-�$���|���]���U�1<��I���]2�N��Սٖ���S%ru�$AcKz��K�:�>�_FXp)/� �KZZ��H��r"�($"�ڮQFa��O���-�I�g�*�A�%�1Hh&��C|��s?���l�`\�}Xn��=� �����3t��i�{S�߃��?�8���U^.g��ge��Rz'_��6��B���ɊY�%%.�j�[���<}�E�7V	��J�R:���QÎ�ӄq����(�$�v�찝[�u��8�d����-Tw�$`�h�%fi��?(�}�|�W]��F47|L�vh��?����TeJ5��J�G���8)w�_���T��ې|iobLدpt[�����]�U���ͭr���ٳ�˷�v�  @ IDAT���� �:��p��a{g��!,�����q�"�+긇��s�F��\6�Mz��jȌq�OE�{��z�	|^��;����^����S<�P}�����5��~��*�ӓ,c^��NQR���2������-b���0�U�V�}�������-�s�e��ʨ�2�e�1D�����H!HؐMq�^��2��@_g`%�C2v܁�_��d�e��@=�D�:>X+��Ҋ���!������2~῀x��u�X�@�+:��Y���!v�C����J���׵��ǜ<}�m��a{1�MB�n�m��qS$+@��jv��b?��F&܇Zg,����y۷��T\�\'�+z۸
�pBwo���J9^j`d]�!�z+�"�8J���7��2Gܵ`�&lC��H�02�P9�Ju�WJ��iGo�dJx|�O����ť+�sFH!酞�'Wg�Ť�G�"(�H�^�,e�㗏(��|02<��-�ρ�m$U9wM<�x߳���9;3E����Z��A�*��	!^��o����lݹ�؅[�]ER̗�17%n���M�\c��9�/l#����F�?��Β��ʃ�롯k|s,��?: 2�9(�h+1CƼ�L.%��2�b�;dX!�2N��DZ�}r�\��wȑȬ����k
F$r�ks�r���4��΢����/����2��&ĪT��,�=*�l���zv� ���x�����ˌ�ི��}f�%fnڋ*ք����^$��(h�!����!�	�H[4؃}$%�-&~v�b�������b,�X>(cD�rEd���+�7����Pgh�� 7�=	�+W_:_^~�*�`�,�=��+�2(i��qfIS���m��8�{���|B�*P�:��UmB���$�u=H��qG��&)�5wp�i�B1S����~|���ÇD�:R�?=L$��`Կ�ն������*;65A=Z���BF��ѣR���B�{��8���!��$;�o����W�Wo�'�0����|v���KsẼ�����<f)��0��x���Dn��qH�0�{q��Ɵ�g�\�U��LL2ܓ�Ҵ�-�+���,�&��QP�b�s�aucN$6�*��%�D�#r����.3� z�^�۸��r|��?(o�vc�
�!��fGe03�.�4�\�`�����)G#��$2�����z�^���怼k�)��3h�ىe�f�:�7�桶}|\�0��Qk���&��2���`����41E$,T��6�y����@Y��}�	d#���r�p�t����p����W�[o0%*�*�ތ��2z�+3�1�8K����.I�	,[�PJDd2�A�M[3�b����A�M#+���@�MS'E�-����g���J���|uU�ӗ��xgc#�7�F��$�˰���/<�i �aV�E6$�E�M�>���׋����U�e0�h��%���I���_��En ���g ���8\�1lѲ��Y,��̎H�u���h%�>����w���r��@F@�5w	�=T�^��/��ꣳ���yT<�� #�/�����s!D^J�	��"_�%���M���+�:��s���e��r����ט�F��	U�خ-���p����8�!�"fe������4�� 6����4��µV�Gw>-�1qk|�1Ĩ�-ڷ���i.m4���>lo�U�������9��L{�:�l0z>~|�0(�x�b�~3�#�?u����{���o]+�}��)���`O{�p5�;��R@e2��|�f:��\�a�bp��&}0"�ĸ8^��������m�'�.��Q���{k|7���||�Y���+����Η��w�}�����!\ơE#��dd���K�H�{ F8�Ctx>N�3MTaTD��������+\��~�T�'Y��G$�Uw
|��t�~����9��.���!�aٶ���m q|�{�
�5����kY��ٿ9@'��f�}������#�8q��4�~�������Ȍ��l�ѮP�Ɏ�]��L�H��2��8��FL6 �[�U\:�>%�:<4�1���X�A@��@��HБh8|\t��x+C3s2!#���x��|�!cRJ0�[_3f&�� v6W�{���*3߆L���(�ӧZ��8b%�n?�Q����3�j	���������Ҽ��r��Vp��0�B�1����럔�1�kw���v��#W�cjf��ch�9��=�<�aؕ!� Q���b9-�7V�>4v���� h�[լ!�]�x�c�a"�_`p����$L���{�����۱p����xG�)帠+~�|O&!3�o�F�P��M7�ŀ0XU�gw����r��M�҅��n�lw�C�=g�}��G2�4�[Yd�;˟c���@g㨜Jl ?lO&8Y�.�FQ�?�%c��ԣ���m�ͤdZY�s�m��?K���*�7 l�2ݥ�>f���j��ƴf!��o`����d�m��4k�̺�l�b�Lg&����d����+E�bm$� 
2!���+)yCT"�!�ʜ�0� e ��H��@@���9ޱT
'R��i��B�2�n�Θ�Z?jF&����ܽ�g̼�2{�k�{��|H��s����	B�)]`��NUG|���v1�3�O"]��pe��q���?���j�{kn:�m/sd���Z�>{�� ��\�ۣ��&-�}D�:�|��P{�s8���;�͒� ˪�!���1*\
��0�XfM�u"ՉC�W�Ie����7��Z2���\:�HX�j�,C�FJn�W6����&�nRl��h��>��sV9}'�w�������'w�#�0"����NPFێ0,qxk�H:��lp����OO�Q����$�Ԩ>2I|/Z����ܒI���X����:;AH�H���0��Ѫ��pK�xl����P�0��H��G(:���D$=�	�A"ۜ1��ߞ͡�?����:$�������Z�oQN�,ޭ1�8�Oh���� �ҜA]iA{!��Xօ��ڲ�/��[�t��r��wG�
R�����Sኇ��H��$�Q���X��<Z�U���Wa	����F����$�����F�f�a��PfГ��q�|�ϑXz&@P�X�m�g��ʬq>\]ŝ��̯��jY ��1tp��#��`�v߾K�1��\�]`����)�������:{�x� fn���wn��l�og;�x�x� OS�*Lh�-���ȤH=fb�۟�$�b��4(m/��\Y�\��bu���`pS��Tw� <`@iQ�Xy���h�my2�,R���Om��Z��}������@i_.K���5f9!f�5Oa��}�U���u�������l�L7<B>�J�t7n2g��VF`��:��Gft~#R97��	�Ma$�\��u�z�,���=70)U�@�(C�sR����b��
^��0�~vAN�'���A����[6��4LB�Vs`Ad�Ȉ+	�aW��S�����"+��٘�������E$�;,W"}!��mr|a?��~�k��I����&�V�|�t`w)ό����N\׹�����Q	<�/�Am�ɱ<i&���'	XD��t+��f�R��F��ա����P1(Of��������,�t�aT	'���5�;]�X�$�}��G[�.�.���ߕ�wn���p�&��EY�����{��l�}ud���i/+��j��Jd��Ѭ��go�v�m\������z�ŭ'���B��)</��ݖ���0�N�x���+��zY����lKص���'��1�!��"� ����%�>V�fΕ�� �k�F�E�{��ZF����Rk�a=wYMD�8Tg:�]�n��W)n��h��{4��ـU0ʊ> �g���9�Ut�cI�|�J%H���N8+�������'T>攪�3o�����1x'Bu	���	��4�>u�Z�(I�ߵ�e��&q<��K�!B�a�o4s��guy�^�H�k��[���"L��TL�F�>`��jyę��'�SR͙���/gs*���mK7�\U�D�~0A���0�):���pU�2	wo���1��pѲ�E�\�3�)e��"�<򉧼{���s�xH+�zQ=�rU��C�H�q.�k��4��9�����v�����{��w�r' ���Q�p�Ct��u84�y��\gq �#�����No��'9 ՙ�E���V �=w�b��XF��6�Z�H[���2g�Z���L����,}�����{��a�����xU�P������nO×�#���أ�^�.}�%��,�QzN,����aƐ��}����A����D�	�����F�`�Ø+hl�ja�(Ke��~����r������e �o;,isp�#pyfeg�#���=Q��!�ӇmC�6K���s��,o��[����i�~���N��GK��g��_���z�j��ʅ�5ADj� ����WG�1l`������`��"U>!MuIЗ��[$~�!|W�I�����;�}.��!�SJqQ�����~����Q�5�☱_d�Y�&r,�n��Ƶ8Q��'����sd<��dF'�ÝZf���8�d�M[G��w����+3`?���#��3Lm������Y3����h��� K��N��Rf��f̸�E��d��҃qOAENcP�w��nb3��=sg�rE�8�/:�$�W��v\�"xn��rNfWc��Ad֠焩C�F0����=g;�z���_�0tvUa*�;�#�c�20$'�ԥ�^��(k�n� G��QOĥ��~R�>�#���2�p�cNQ���[�,K���a�#$��2�7�Y�l@�x̢)�qUݽ��؈S�� ����xX�
n���SZ�f�1�S�}��UԜӨ������!��$���F�]�1җL2A,I��&�y*�a�3��JO�#ɰd��Y�Ho�H�h�6���fQH����8'��\��6�l�����\�_�gm�*^2���s�eei�ܽ��vU,�X�7Y�9������1M��p�&�ߣ,ٌR.���mmt��yH���x&�8N&E�4�;����L֯~;� ?���Y�=�fg���M�;��o#ԇ3�1;�^1^�"���<ak Q�i�iB��|mJ��FL@@H��2�RF�)��CkuS�Y���ø��R���sы'��Rꠞ��L��m���2&�Xi��e= �5�I��������IЙ#���g�x�� #"�%�.���/'�y�$���C8Q�7����_�������0��`��+�W^�`�.�|�!��p�қ��Ke�s3e�pAz`{�p-��ہ�	��Pŵu�i'R�� 4�O�`
I"���D���>sF���x,��հ_LC֗)m��07Y��.��!l�.5���^� (C��,�Ʌ5b>�gm��:îMf�����>Blc������-yo���4�af=��g���G��+�xn	+t��I]�ܯ��s.@�I��5o��֟O}ۆN	7�*���;�cX���דvtʅ�s�Dҩ�s��ֹ��G�}QR<54��e�@]{w���3�l?�QzGMzBn{0/���Agf��MY��$�cV�6�8�N����R+ �"�������Lg�`mX����.NS��3+��D��T�y�𥍱N��ɦ8��lL#lQ�d�|6璫�_C=�O�;�"�cu�q����?�}"c��5 s�ؼ]�nb_����CJD�>�����YcÓe�m�|V�?�}��q��}�,��1�ofԎR�^8�s�B��G_h�Qŏ�H�� �80�Wq���5����F�B�s�O?�Fw!t�d�Q��Z��>�
��[��]�5��{�c�1	�o�;�3c�:��O�^l���s{9�<�N��jj{!AQXq����zt�
K��;o�U���~�����g�1��j�J#
c��w	������L����T z1�pԊ쵥��[����EWǛZ �Op���Id<��`\��Ն�4�
�l�Q���98�����3�C�H/a��&��G�&$�@ ]z��d� c �3b"Z`r0�|���( �S�h�PTwf�_��_BR K��x�?�m���H����t F�'Z�}`EbtD��a�8����~�,mܡ\\�Q,>f)bk����E"���%�w�y�%cڈ�u#e�i&6�����"ȹf˵8�ܱ�hi�yͶ	/�k��I�x��l�Y�D%'_9&YR�鉱�:��AF�D0���PH`f1}�u���VOY%�f,q�j����,���*���s=�Ƚ�D��PqR�r;�����8��+s��#+��k�U����d(�٥�k˻S7����
�	�_��_ӫζ"/��cZ=]�#�<p>����πH,��[������$Ta�&6���	n.�"_ 3�Z�ƱG2y(�Y�٬�Z��wz\:�y&�"�����3Y��W�O�Ђ���c�Ch��u��PlC�|���GfEsS�:�DN�x�;�cM�����n���RUy��Y<�q��@��J��Y|��h�W3b� �.�,��%d>�j3��!�]:l�8�t|�(5�F���㋆F��5U��N�ϣOR1��m��7�r/�d�Vi�NZ��F��zm���A�2��P̠�_q��`t�r�USC��!l�����K/�l���Sw	��@��|����1��pS��13�[���t�^g/��u�ph���)�N҈�?}98x)�Y�Ӻ�sٗ;�X�e�y?����&��t�r�!Xd�HݏK�ѕ�9c��k�P ��H}�7��w �"}�F[jap�w��8�c�B� w��8K��������%�-"�Uw/v��Y�(�S���U������Dx��i� ���k:�%&nl�� �cV|�;6�9xNjD}Dp\��f�����NN��3���c�E6i߱�g��l w�ʐ�29yd �׭�ɀ��%��`�9{W	@�*�1�U�Ð�x5ʃ1�'�)�D}J�!�
w���,� ��[�C[{H!��Q���*�<�4���o����?���k���{w��P��wF��h��2�/�a+f[��ѣ8hg����8Ssn���>\��
��6^`Qq4������x���|)?��UNڒW'9b��g����mw%�'�2:�r-3~t�����s.��ʀM_�"ö�@~C��| qoo`�hc��".�D����.�PF�!� ���V�1�|1C�N�X�E�<
ۇ3��J&�qi|�0�k{�A��P�:��|�x'�ǆsOXADμ��F�H��o��$�8QJ�2��m���]�)u�όΦ�*m��،��)�A�1<���K�$l��>�!����Gwr61Bx�z�S����\!r~)�PG�ΐ��j�=��Jд�&XI�H	$��(��/�O�`��qnЂ�x���)�U�kKv������[Ve�7ơ��
�O����Ku�$�b?��ƌ3΁+��3Efo��}�{���}\�y� u�9+�n�w���?�8k����%��R�g�34����=��{]%t��}ݕ��R�)�*���tRB�c`���L�Ν�+R�)�JB�8Jg���2WBD���,��w�$t�y�3�4uѬ;��*#3���I����Tڤ?�B�4f�:����k]ά��a����H�����5�"'��$�.桄��ϹoJ����������(D��h���������(�x�k$e��۳���3��(�?��*�0��
������V=��(�D�y&���3��X�d$�O$*f�vl�f��
�[$�`8J+ҡ����0��`��;v�"5�)©~f ��i�Y�l4[孷/`�a+1 ���Yp��h�D{�����1KL�qp����-k���r��a��)�r���0k~
��&� D����&:��;�������\���/t���T�[fW^�A���E�&(�,'��VHP�`s� ݸ���&+5i�����"��X�p,ESjat�ܤ�}��# k��_T.�h�94RJJ��{�X����O��B�2�V`#�}a:<	C}	f�R�<R��Lؾ� $l�r	���+Jk	�q�����,�Uk�ђ(�m���iK,�y���Q���ϊѮ��,(��ؒ�Q���jI�&�s������ӻ�]$�%kQ�p��u��M��<�$\���J\?���T��_��CD�U�l��p�wY���YZ��Q%ҳTiİ ����so���t�}����ݲzu����!ۄY~
�тn��[?���z��;���wě�g�tHHǜ������i';�uԀ��`Dg��	D�T_�d��%*f������[�U�h7�x~������b���;��%ey�4���-�����9^1Ȩ�Vc$T�~"�D�`�)ID��Iâ��g`|��a��6���;��Y�:(�f���P��(V�cdRLיJ)�G���|�����G���k��s۪h�����	�
p$���t/� F�ρ�@B9)3�jV��:��6Y����2 Q�Bo�r&h��9Y��Cl6�f@��_��Q2C��݇$���O��XNJ6>�?#��fD�N������XH�L�a\�;�<~���\��w��ڈCM0���x�'�l����=Cq|�xs�"��/��KMC,��6�����F�������z
��<q�:��>�.��߄V�xW��:9=\~���h�8���~$W="�OY�4V�bDq��UW�Go �C0���!rUn�ӋQ�t̶���wz8%��e���7�a�bEk�Ved�� kL��Op9���H�{��P�y�M��C[� �ZO?��k��l[!��lk���ry�yh��;�c������Jq��!R"�ܫ?��'Dzo�>����ו�z�s@�5��@2�7J� KsD]�#�M� ��;k,JW�lI�J����$a��e�&�[�;K�&g�˾/��r#~��X�pU��]��W�_mX8	�����c�=�?�����lNR2����>�%� ��f���a��W�I��`��gzK��w����~2�4E 'T���,s�܁6�>a� �`���Cj%;�kl����w���$o݉�"l�	z��>�e�z^M���)mP<��aw�*�q4����'�q�-��[�"W�o'bS ��	l ����j�f�~���uu�F(�C��/����\�ܬ�r^g�0���T����+o�O�}l��0t��O�oq?�H"*���o�Q'l����Q������7!�	粚I/X�q�}������F� 7�a�A��D�-�	���=������纟Af{��{��@,�����Q��������Fo�~86؞bF�.h�����^Mq	��-ɖe�@�#�J�M8�6g:^z���������+�R��`���x� ����[sz�<9"<`]�L�3�n�q��+UH���b�*�y�M,Y7�4Ȁ�����0rS&$��S�l%����RQ����,�4���m-�8����b,��}�`
>KY~/5U�+����|�)��+�r�$��6ʰ(�qM) �~��v{f���L#p�]m��ey��g��(�u��PS>��
bq�$e�;ƚq�|fm�K��,C���>)H�Q�)��+����dx��,Vk����1{���㬕�i�z�\���oSD��1�&:.�d���3�H��9b'3 �m�<u��&_.+��<�6�#�p��@����Χ��K0F�&NK���5�^����,����.:�O���F2v���Z����Ѝ�C�;p9c�#�����02
q��x�%}:@�5���a�2�\��7��*����PUg|�)h��P-Kh �6�JC��AxP�3���a���'�䀝��y��C�g8Z��#f���Yo����6Nj7���h�����k��;;�zH:l?6))�j��jkԎ�QH)Ü_��>��A��v����8��3��C�x���eTCK�D���Ý PEɋ����`���A���Ҽ���e���ѮC����Y��
cdr<\�I#mΨzo*�dyf0gT�E;u�VJ"Ds8EA���m��v��`�-&���P0/a�H�G��~��cʛn/"E��Ӿk�x��0��&u�om@�����a��x�\�Oi�t��Q���|	P$SՖe c�F�����33�
�c���?��}�/E��F$~vz��cmv�Q]��S]fcu������5���Đ8�ַyOQ�D���7`v�6PQ�qfa�K�CTf�5'�j�W ����AA,E�m�i�Khw?��k�&;��?��Ƌ�X���� L0�o�RQ� �I� �8��$q��m��a~"is&�#���߀�PD�R="�!�N��fY��w4�2�㜀�D۬#:b��ɉL�����?�#f	��Jc�,=�H���@�����n��ĺ>��I�7��!���IT2%.Z�\
��2	&��~>����	�@ے@���)T�f��
���G\�.��J�Al��̕I��F��!��ݍ�8�i/��|@z� ,����E�ZU(w:Z���y�l�2e��/�e1�М����$�ʬS-�^l��i0��2�H)(KJf`-�ٺ�.a/�z�d��՝`t�,��w0`�%�}t	�=4��O�����:v6��~�E�I
��k�J�jϩ���i��@�������_�s���
��@���߻�֏..R�`�x㍷ʣ{��0�,g	乽?\��l����ޝG�x�3�����Y�9ö�͟���ًd�,̟§b�^�]z��Xz5\uǬ��~���	�!����'oZ�Q+6��)�Mf�+�a�v�g�Y�N�
cc��;H�ۨ?�>6>ɻcAl�������at��o�k�qu8�o��� �q��؁)�#NLP3�����>ڶI S�cס.�ì����E�@��A�I�"T$�3���@H���(W����;����;��+g_!��q����n�Rw�s���A��D��l�.�4<$�����G1z�m���jx�Ё������.�d$\Qӕۚ���\�4�.󁂈�-���*�,�c�v�X��Nv��<�o��@�BY&-S8;������ƹ4��9I��с��|2�?ht�,�W�iV)�*���	�w��F�_��e=ɜ(Q��*�{ͻ�)�v�Z���@�Ӭ��$s>Q��V�{p`�/㮥��;L�J00JT"r51��;��AlkH�rsˣN�>"��활ƻXܹÞ�o��Q���O�YbM����F�9h3��E���N�C�x�h���!�uY�cǶ����We�ӗ_�2��b ځ��n���k+����!��������V�1;��+qo��F��-���֣29>���k��p���Nh�����~�����>a�O-�*w���4A�S���0�c�e�52P�pb�I��;����z!��P�9#����Ç j�d����G�e�L&��=H�Ⱥ�c���q��\T��]�
j$-gњ�.I=�����x���O;�c�@?� e�߇�������9]��������q<D�A�]~v����q�"�A��P�J�HA�ۨ�Ee��hZ�,�T�	q�l���ڀ�viN�tu��Eh�Sf�<l���em�]�G=��gBv!c�%.��]%4��6���g�~0	�����vr���ͳ���K��oIrJK�͵�K�Ƽ27��j�Ax7ꃐ�|�{��x6���4�� �e��\��yr��e+�N����� �k��w��|_���z
l%x!I�g�w�r0fr�S��~6�x@e������ŗ��Oo�*��>f 6�`�\o��Џ �k�;;�����s3����Y�aY�𻜕A�u�C�#j�n��� ��C��Q8�(�&ݵ7�-}���I�����Mf��7qTi�X�&���p߇"�
�B;�t|d�駌q��a�����V�: 0�~�6��xPF���W��l�Xd�q�1m%��#���$�\��= ����NJ�z�=����%��}�8;��������1�����=4]~���Ar �侖�a�f���D4@h���2��2q�X����ՍCʥM�>�Iy���ڙY��%6)��KS u#�G�K �/猪�b9�>nuI2��Y�Y��kt��Y~@I� �Ku0�<�%Ղpf����^7j��h˰>0������{`��m� 5J"St��1E � >�X�&�K܎3tPjS`̖dDq!���Ȍ���AY��K����18a~ۖ�@h�G�B]2	��O2ǫ���$ÊD��d+-K��DNO�2�#Ƒjy�Y� >$]WQF�y�H%�
tb�4�;9	a��c�o�b�&�N�5�@�;�j��W(��a�m kuy�,-�K���e�r�H������-����sJ�k�fO/8��|D��q��Ә�}�5fW�Fi���K9��+��T�����&���r���F�R+b� �DC� ��T��ɜ�bx��h��F=g�}WR�A��+6�zl�l��@�"aGO�"b�ؾ��	~�a�d	�F"BǬ������*C��M�M#�L]�1*r�-� �>m٣.#'���MQ� �L����Pۨ�(E�5��1Lj� ;n.Z�<Q"$�t��ըy ��܌�`Ch-������2<{��A2HC+��*�ΰ9��R��a{�� 
	�*1vY1�	�m��H���`���?��r�!1H�]t������ROw��a�ΒJT^����S��1�\��.a2 �C��Ūݨ�q���J�Ö�{PM1���c- F��Dˋ�9T9�v!��oa���W�  �b�]ڌ]�T�L�*�`��+��[��$Y���%sS�@P��v����ב�|��;��Zj��h�h��ؐ;Rc���n))�%��w������K���$+~�;,w8d`S������\��Y����Q��_�$�c�vyO9�9Ό%�~�a��.�3���<�Y�1��".�Y�h�3�@H�,�����5qy�s�Ft����G9�lugy�m�0����27��&!ɷ8�h��"3*zsހk��v�=@��!�+ei��cX�ȳ��1���Ѓ8���g84��� ����|x����-럄3L���1"����
E��bhuxz����!gP��Օցz7G�l`�nV[�>�Xf�GzYY�O�Ē|&@P�$��)��t���@�������ѕ�(�(�qer[�K����rH{9{���o�L_�f��H��sc��Q�&G�g/8��G	�v���f0�2��F?b,dX���y �4�����:��"h}O��`��(l��`8At d$����2�5b��8�'�{m�
�]�{̡HƧt�ML�栽LF�o�ZY�߶��M��CҐ~�.�<�.x-e�i����HS� X0yDA�`��L����,�q^�`gZ�t�8�H�T����G�l�wb��j�p�@[���D����-�g��:��ͤ*� 8pH<��#�!���B��mo�p�o��{:o�.7��P�Q��SZ�a��(�S�4AzQ�9�P��Ė�_�?W���o�xθ����l�:0�����,�x^r.��7���ߡD��Ǩq6Y�8~�4�M�p���|��c0����,tn����Ǭp#�p*���/��V.\Da×�84�=^����2��2�?��[_����b�.+������/�f�ى#'GX����N����w��D;Ĵ�*�Y~�:�;�F5w��!;���8 h�b��u|�gUfN�
�Ħ!ˈ]8��tl{��NY�`x�@"8C�.r@��}f��s���6��L͕ǟ�(�ΜG"���?��΍dV�@|p�QY��l���i[������P���,�>��r��W���NNFUY)c�~<�8�S"�+���>"d��2�4�i�È�k�'�@D���`sC1�Yb6G����(\�Pl���h)����&� dP��#@
�Sx��{.g��b�Wˉ�����p/��$�$
�ޓ8�m^�m�2�G�j�����}~���
���і�c��S*��<�O#���A��mɏ����h;���$r?��#	K���1	�\m�k�Ⱦ�Q��ea��]��!����*����M��K�>���v�x��$�B����+�|Y�C��`H0�P� ��Ia@�[�I&ރGi�}RR�d-���+��hk��8���77��}bd��_��elGe��Y������v�����1�1�|R�_z��Y�B��!����J�cT�}a�Cvge���C�%�����ʷ�d�f�<�cEG�-{�h4!����2�� AJ���j�揕�J��� ��=�^�G/2s��i�4ڃ���L��<�.t�Ls��0ƶ�;������'�
������c$��K���Y]����(C�`�١��_{���ޜ8S>.�)��F7�v���K�J[�7�6��0PN{�b�<"@jK��Gdu�`��2I�d#0��}�`&��i�*0�^� ��8�n�����ݨ��$gA�P}J��(�������Q��w�8�K��#N�*/}��^9��<�D��بخe܀%�Ȋe�Y:79��f�<�H*QH�<a%n�EȤ��'�%��ǳX���Hq��a7H�"������-����R��)"����B"�}���l����C�=�>�������s5T���oG�˷:}��3�~yv�(/�M��-�AX�(|�G���Qsl�ua����4a�AbL�&T�D�cs��`0�8g��l��	F��J[e�t���OF��o�;�w��}g�RB�y�~�]�b��a��}�,�*� 1`�t�^���z��w��>�y��w��W�#�9������!^:e�귡���Ǭ�l�Y��k��w=k�S��C��k�v{���'`GE"BH V��8@�N9q�9�9H� !��Q�۱�힪�����i�k�5������D���������p��u_�����_��ީ���G	�럾�t�z�FS���Y��ͨ|��Fu���B�w>�����Z�ܹ����
+�㔊����V~�U���o.����VI�B��?���̇��?�xy���?/��یv>A;�?i��������������#�:��ɏ�>�Lȇ�s?F���-���������]���:��'�]~��ǵQ����	�_(���7��6R���]���fT����������E4���wd�;r��%^�(�����>hXTN��_�|�����_>�����Me���r=�:��\��6���'MW����'���.�ꤨ���x�����h�?�5�[�s���q'|=}t�򝯿z��W~%����hC���
��72����V��$5	'a��G�M��٭l ;@Ŀ%j�k+�ji����V<��^y���8K�J��z���꣧���p�S�m�̏ꨡ�4�NqK��Hd($6��$hJ�t��螷���Kp�\柢��%�u�ݫϺʷ� l�jFq7�L��5����oh%�H�M��]��l�AE�b֮�3/&�Wm����86�q�K ՛��cWFb���%?�@�O�35��1Vure�.j��P�K	޳��A����8�/}�s[�b��Œ�F>_nmÃ;�
����/�KE��py�ײ?��o]~�'���,�U�~��-7�5Vz���������@̬փ�ct�D�?�sy%��a���<9����ˣj��N?z�����Qȝ����_�T��-�U!ُ��#ҫm8{�q�7��_���0��Ƿ/�����T��g��o�H�����K�5�����z?Z4��݋)\���k��^~����)�*ٓ��=�  @ IDAT������Dȟ�{��?���<��Ƥ	���|�s�y��a���7�j��A��D�������߿���)N��'��6��f��Wn-�۫�lK~��D�>��^zry���{�"��/�336���^C�O5�z����k����>�V��������|�����;k�5K�c��I�=���q���1�3�ޙ��)o��o��SJbJ�M��eû5�̋%�}>
�����C�b����>2�[�#����Ez�:�l�%08!�w�na4;A�_J��6�kF���
b r��N��ζԎ�؋�R����`ORj�\������]��CgI5����"ҘҳF��伹kU$�1X��z8��[�^����ڹ�4:_1y��\ƆͨM���yfd��(n:�A�ܶ�#:�ǻ�(����jX�;�݁�k��J� �ky�w������˟��^~��ou IS)ˇ)�˟��勿��u��˗���?����~y��o^>]"�-r����)��eg뿊��-��T̋v�5��aӗ�>*�RBNn�\�l3��N�)����LC�X_>��^^��ޤ�^J,�x)cb�全�9�6��z���ہ5�>yx�D�|��^�}�Q�Z��ƛ����g�>�YIQ����	�P��@�T��G��ҕ�p�
������z�{�A��W
��O>*���7�F-�W�;y���x���ů�R����o~�%,�y�8���Sc�����|��fm��F9�؛�w�j�3
�Ey�'�;۠i҇O������v�>�<�nV�9nj��W;����0%x�����T���	��!YYr����\�h���0�����?���'`�ܟy���(�
��Hm<��R�ކۮ�Nє�G�L&���M4C�y�jf�♽���:9����������f�ז�!lw�0�[�qU�mo�C�,0���D��ވ^���|�b��S�]g�aL��oW��Ul࢒Eu��E�uFS�&7��Z:��|����8����k~��K5F7ѣ�!�'{qNhj�5���?��*�u������2��/������o�ۗ�>�����j��?�<�=��[���G�(����+���V>����75�*=��"�V�=l��3�����^��w�n! .�!��/��Ǘ�{� ��F�?���j���D�AK���po�~ء����e��k��:����a�%�%?)��~�y��ۗg����u��g?�5����i��)��%)�x��ˏRҵ��|�~	��G�����Uz�|���|�"�����~㽆���^CX8�r�z܋U�z�+�o~�6[��Ϟ�l���[���E������<-'�{z�{�w��6����a@!���۽h�IIė�o5DH���[E.�Ixڂ�[�����<���S�ߟ|+��������K��۳s�e\���&#,������͌˯����]��^��M7>�c���=oz؛�ͪ��fP|�f��E'�=��b\�&���a�|�bw/!�x6�&�9�-�Nզ��_e��~u���mb;S��KYΔ��yX��̗R���F�?	m�����O�BY��__�T��tl�8b�R��L�����L����qn��7�[���:�	{�`�2\�E�p?���4g#��o9{A������E/�!|��A�<4�A�C�.SE�X��6V����r�[F<��Ű�E!��"<21a�0�{M�}�/\��/�RQ��M�ݹ|�U}��޼���%,���/���ry����/��=�t�$�z�Η��w��������a���.����s�>�|���撋^y����^���?Ӻ�� _������{�7���\��<ާ����W������������ƿ��7-���;�����~��'�w.���rO/�?�?4^��_�W�b{p���߽����������x��˗��_)�y����7/������o]~���zk�x�ʗ߻����������_�H�_�����$�{����߾��������������o��������_����ry���]�|��i�ͷ>�L�.~�]~����k���v�~������ft~x����?��Ϳ�_���O���w��.�o����������w��������Z������o��%Xz��W�zy��\��?������.���K�?�k�|�Ǘ�������uy�"�w;�~��z��w?|��y��w.���\G���_>��_lE�Z���ˣֵ<k��ƛ���7~����f�~��˛MyNp2Pv�>��fW�%�9C��y^���� ����� R�"��];%�d�y7�"��ϔ7{����t����y5�`Կ��-���)��+��"����?���Q*��-�V�n�6��!7u�59���h��GST:Ǹ��uR��C�NF(E�ٚ�pڵu$N�b<�b.D����o�;��4����=1�UKַ�>|bD{�,jP�z�*R�.�E7�f@��E�cL��!ߏ]���-��0��g�2����M�)��zɈ3��+_�By��n���R��_Z�z�NS�_�W����у϶�plK>���͗��p7cR������1�~3�M��_�[���:틭B�S����._��M'��P핒r�����ߺ�o�7������?����Hk"��G��e���7
͋6�/9��۝>��؛�z�ꝿ{���_�k�F��Mi������O?�q��f
��y�����+�������������_��G��«_���q��O���lY���\~�W�P��G����7/�����˓,����L�����巚z��z����<�I���/\~�3/V�����?�qxr���}�5�[7���7���)Oo������{����ӆ�7�����w~囗���ӄ����O/���'%2[�����?�Z��}'6�j
�[�����/_�'	�WB\���x��F�>��/nz�E���6=z�%�.	�;E9�r�-)�\���KT��`���L ���<��!�9�jOIk[MS�wL/uQ�)Q�li������_l�F�%��A�68��zN랍v(��ER)�fo�J^��";V2�G2Z�bLA]�?��E��Չ�y��y��Y8Sp��j�ڔ�<�Vu$�iy7�n��wwPt���6��w� ����T����%zEuD��,�c�������}	����h�A�\��,����0��9�����^��h�R�o�����r�}�N�%�Y�������ċ����o�������������.����˽׿p�տ����;h䭷�Շe柽z�����2� dϢD>�o����ӂ���֡?���jz�aY���y����~�W/����Oʸg��J�����_�+��_�\��2}���KZ~|��7��d�R�JV�Ny���}����ʵ��靯f?޸����߽��ۗ�F<*|/ur��;o�g���������^�����|�O~w9��o�sy�d�O:|��%o���Q����zg0�����]�����	��S_i��Q���>��WaWN�w8�j������g߾<��'�Ͽ�TgD�:�̷{��[�y5�kH�����y姽}����NÏBK+K%����b����ھ��_~�.M����?����ۗ�~��E?n���EX�M�YA�"S�	Q��A9�2/C�yp�5�*����p�沇�0����j5�d��"�7YqG�����D��)y	��Kmp�N2+��M�~������ TIIY���bZ7@�M�>i�����Ĝ�ȌDt]���@QTpDϚ���)���?�7��Dֺ�CtCuE�$dC�����S0o{VD��NC4�A$~g�axMF���j���c��\��E���h�Bd��#�P7:ș��������"�L�xU"7�{Ql���^�3�V4gQ;��[�������O�������\~���?���+�*���ǽ+�N;�x�˗��A�,45Y�{%���4j��	�GvDbp��${Ԣ�/�����>��E��~9�ݹ���~u�~��5�{=�}9!gtl����L��~�-���/����������j���������Á*w�+���f ��b�ag���|����ԓ�<�g��O��O5�Qx�s���Y'1ŝ���׶�{alS3��:�RVުA�R�)_�Mi}T��7��X�vUV�"?��ݒ�	l?7,�f�}���>J��G�iS��}��������N}T4�5�6��c&A����je�Chm��BQw�s?%�F	�;��;��>�ٮ���(E��I�(����م�S�zF��k8�����j8��
�f ZsU� �n)����!)O8^ԯY�](���}�/���ɣwQ�͐_�hE�TP.e�0|-�L��'*%Gpb�,r�t��[1�J�k�k/ի��JTG�"�FZy���5K�.	Lb���$�)��$�!�1~]��[�~�Y��l#d���"��V�97�j�q�Q*<�!�Ѩ�_�͠���n]���W�U�� ��=���[͋���t�׼�0���A�]"�q���<����g���f"��6b<y�}�Hu��,9���$[�q��~���^����;��_���'t����氫��|�AS���Q˂	���&|�+�Yf��9��~q����wZT%YTD�Rn���g^+Ri&��S�*���ʯ,�jna�R3&o4]k\�Z�~�"�/���W��Y9���'y�%՟$�Z��Ճ_�������w��D:\´Э8��E��f">l������^J��˵��~�����阔"�(�,^'Iun�k��`d?yڢ���������h�/Lq��֧[)jf#��H}��7۷��a������R:��^K����&�父#�A�X%�� ��.�M�6V�d���Ă�eX?n{ӑ)=`�l�ӆH�i�gi��sWfS���S�������=CQM�����y��;d��7K�c#Sj��B�xy��ц&B7hS���Ӕv�Q���W�j̼0��(YhUS�m,��R��epk6�W��V�w���O3��%���qM?x��6�~
�U��f��c�~�EB���
����;"Ng\w7~j�9�pc�j%8�7$A'Q'�N0�Sd$k�I؝pѫ�~ZH�F�'oҽ��G?��z���S3e�d	�G���&��?�����>i�� �{��{�_�;b��_�ɰ��K����qF���\���"�W�I8}��)x�x��\��=k�"�Kl-���E�2E�)g���~�з5,d}?5���o��Ol��z?�	=��7~����(����
��d?[�I��~�����Q3��3�3��=���_{}[�_KIysKs�x��A'�;�6|=jx";|s�	��� ن�Ȣ��a����^���?z�{��7��q�'Q6Z�<>�;�R��y^�A+Q	����N�	�D�׉�T�FP-����3a��׍B���CS��M]�\�b�s)�y�An󪔽��}���Q4��t���[�v�l�]ЭMO��q�пڪ\� ���M�d��ﭼs}R�:̘����}��ڮ�,�u��X�e���f���sL�R���Ё�=9��P��EK�Gݬ����*08���K��(�!�9Ȩ�6�q�ڒuw"���8:c�'��';�Sy��*�g�q-�<z�f���y-l�jҢu5{��kͫ?��CP����_?�Ƙ�9���خ�)�����aVRg��|�
���1���-W�ߎG������I��V�b��~���٘^|Tx�^�K��0o��{Ǧ����~�i^d0>ՉV�"��Ay�b	�ڹ����,�9�W��?yn�m	���w3\�;�B��&�w2B�E�:�	��hT� �_�|li�K��l�2q+���1���t۽�V^��!����0P�Z�f�֔<�NՒ}s{	ie��3&J s�n��Y�{��o(o��~M˙6�ᴿ�`���X������v��2�ӿ%ή
����ޢ�E#�V]�0<�*r
ohp���.�O�����9׎��8m,���RΑ�1~ƫ�Ч��K�q����Y�_4r1��P����QS<ȣ���΄ƻ6yuLV���a�]�w�΢��ͳKv%<��6B&�e��o��Ϲ8,߁u��ϟ�A8YcE�p>|���};���g�G;e9׾V^��>��a@
e9�?e0��1��`x����<����{�|�X˺w�F���M%&�5���;Ü;y)�Rv�w^1oY�#;�P6��ԩ<d�����5��1���SXc����Nr~PR.:��hKs��m�h��I��VC��-�ݎ�Ƿ��yj�@r�&�3�la��Z�D`3����z�����d'@�ޏ���J'A;!h��-�e�^o-��X�F������͌"��Mт�A���~0�&ܾݐ=�,�j��`�ۋ��_Z.�=��ɳ���k)�z���b����A�*��ys�S�ㅰGh�9�S1�^C@᣼���7�Ӫ���ϐ�L����T��{��I��1��:W����&ԯ�)�B�3��"d��h�0�G��G�������<ܕ����Hp밟�<�+�G�ɿѤ���$�xV���tϜ��8ph��L**�U�E"o[����xPR0�"��%�G�9��Q��5=[y��n"����Ilqy��͒��?{jG5.�y�v�1�K�ְ��c��x�s ��N���u5���M��A��peܢ�����}%~�1���W��Na~G�9���a
n����d!Jh�f��w�l6��y�ba��f���0.��PR��^n����^8���-�u��I��i6�7�+�2^��=\���������|ae���风�{���j�6��n�+^�&�:	7)�;�	�Q�&^<(����R�O]e3�`�"<ź3�$,�a�-�~�u2¼񎿟�brش���Kx��C�����:��~�y'�t����-�(���m�~�d�c�����/��w�ٳ��9�61����/<K�z~"��H��Ԫ�[EJ����HC�*1?�Rqm�X��^>"ػYY�S7FBW����I8���#�Q$�䩺�t�$a �\��U�Z�XS��1��&��w}5��̵]3�k�۝���,�F�rfZ�y���0�W78h-�w�6�q��[�1:���2~�k���`�^hof�,(�X��!8�"���km$Ѻ�����iZC��%�;ZJ�V^�Tk��_�2~k_OQ1G!dh�v9ǻ7�&4�9!��GMI6]x/B7:	Q�I����BT��~c]���5���	T;�* �z�a��V>"�Pl�qk�imP��P��,磶�J�j��H�>6L�d�-���,�YX��Ӭ��4�m�񽞙�x���w<��jIF�/�+�+S�Ic�{�')�)'	�W_k/	�2.����@"Q��2�/e�	�S�>ns�ĕ��-4�8?V�8Bt�T�#�Ǘ��O�Lh(�M�yA�CgoX݈��0	˶��?~Ѹ�8s��)�q����wD�2�阂�c����ED���E����a6��
�����{�/��#�E=*4�6�Y哈�xr�=$��͓�����o�/�/x�"��"�gB�ŜT^�SEIj6�]�)��o���
"�~��c!���xa]�Ff�ӁG�=��:�ʲ�t�b3�����#rG�<�w�X\>V���^�ߓ�"�$7ԕ�x1xf��C.O&��mk�3���.9x1$������Yы!�3Ul&�4�����K.b��2�W>mȑ7Iѷ�-�c�:^!d�Hv�{�~�GXF�H��8���T�h�/�l��5�����7�:��F:		;��)��� 	>�I�B���e��W�"��J�"3TBl�3pPF'8ukB��*�@\�`��:�t8����L�L���2�x�o�<��?��':�z̌�ˎ��@P��DT���܃'��9ª��W�}���6/�޻�E�e���������V��p���ڧ�7e����c�waxE��#w����zj�,	���aK�w�E����Z������#SNt"E�T��9��w��nDA������6t�8�x\��y���et�{x�]>K.�&�+X�s"C��P�kDkr2.���~o�%@%#�M8��L�Nh�")9>�%�r������K?����ށ����F�zyQ�e�pw1`գ{Os8�������D)���{�f�	���j `+�t%��1�0e����D�Al�0�?W� kL%3[9�,����$����}}�n���Q�"���D�8�7u:��s���H��O�\���>� �['��j꾶=��m겷�\��`9\q5m�=�S#�y��:O���j~(p~��6)�B}��#�JN����2Z�V�}��U�������cl7m�N�Bk���co�rf<����U�n`_ٟ����"��m\����b��P�a8�C5y���P}Cƈ��½��/:�����Տ����юq��E~j5��������<9��ر
&�R�DwDC��AS{��zF���|�[�tQt�͹ʁbmV�fq���)�P��i�T$���t��0Σzt������[o�DŢ��S��J�ɗa^O���c���s�n\���Ю~��NZ:ɀYos��/m�p�"v&cV�搣��Q��./l"\,Ѽ�(_�}G�O9X� >¿&�k�����yp2���/aB+��ˍ�Ow�j!��� c,F��f
��G=���.�q��ڧ��8�ة2�8:פ�Ԡ�Q�-�E�ڝ���A9�����+b�u@t?�aT�ρ��H��)����SJTe���1����h�2�f����O�(u�>+[��	��eMa�c�a�^��u��;�=�J�ӱj.0��!Jv���;7�s�3���ӝ�,9�й��n��e���q��S%=�qT%���^��E9(�`��ͥ_�n�"�m��*���ъ9�0PՈ$�m����!nǈW���pv�(�v������6X46�%?">���hh�a�T���j����dvy��|�W<N��+��͢��!Cbvp�T >3.c:�Z�Ƃ~w*�_7k@�}`�"[���Np�ԞBG�;��6��j�"�i��W� q��xLV8�BO�jnAH@�6t�\=���DDD e�:�q �	,���8I~���Gom20�F��N`c��o$)��9*U��p�
���c8tf�#�����.^��D�BX�,s�p'`���A�9p�!�Ť��$��y?�e��~�����ϩ��1<�ɨ�b}W!����e������enmBĽ��D�c>�4��+�kS[�*:x���bS����d�6�����i؅���0����y�Z=��Z���yj�<<�i9�Gr+)��֦�_n����k�0\�
\V�Z���~�����@|��Q(�[_�=Ù����aĕ?��ڋ�d�e�����0ڏQr�K�w���Qy4K��P��9F�h�Q�%B��V��D�v��6,����9�����Q6�wWۓ�J1���"@��eAO}����P0�Or��ŋ���[I�ڃ<���_o�Ke�5���2Qȹ	�3�@,�.x��<L�T��-���s�j��sw?�Oi "\����{���%�V3�q�Ү�kbZ�yի�"�~��,�}�Fu�pLC+����QDJ��K6�T�)p�1̞?j�0�E7����&H㡡S�����/�î�$�H�7	�~��Z��uA36F�������\p��84�w��m�EW��N�pGmt�3�X[Y����[�A�"�ֺ0��;��wKhڬ��x��/�u�gW$JO���βh}S����g�?g`��t#o7y�=�L�'�n��̉t��)*ZD�)>g1O�Cq<�!��D��K`�-�q:��M���'B�x�����tj.^t���1鞺�`��X;E�����Z2���=̂�6��1��l���KĎ������]ҧ6��ý�\q0�]6��8���pc<l�m�X�)���8%��$�V����WI��S�_������<�	,E:�!�$Q�z]'�}E�� ?%请5��(��^��ʚ=��h-u�����3*du�;ψ}��3a��X�x�Kd�������ǰhC�)�*��/^�W}MȪW;�%�2,hH��z	��Z\���[�w���H��R��2�A3���h�A;��»�9��:jQ��nC֓BZiQS�	�ffD^�f�ɪT��;n
������p;�
{n�J�E��
�j8�aH�p-B}ڔ�Ȅ��k�2� 5ݍVͺ��u?f��X���������&�p�j����U*O��,���S�v�<D�:2u��v;#^��{OF��`(�@n0�.Y���k�Iy�<ϋ�*���J�*����󖙜�j��
�R�5[@>�N=L0��>J��C�'�]R���1t���9'P1�qͭ��[�d�����az?����u�Џv�ܬQ�#�G �B��f�*�w�����T�vneO;7�-���!��>�>�����*����%�a5�,�0�{%��	�� �ٳ���Ϛ�3��$S��8�vE+1$b�9�/O�w��	Ν]�_��_�=�����H��ZU��v�7O&��.���7SZ3���3ޤ���R��Nv��W���>�բO4�\?�`�=� �����g𐠢1��������ג�W��:�*�E�=�� eF��p�V��d�H�Sr��C����rR��F*3d��f���D����ՙ�Br�:2J9��)Y���2����/����&3ڰ��K�>��M������#�L�k��$��3S�h��^��Ր|ӟ�1�qhXǰt1�V[�{�A'��D�%\�6����Y��8�hx1F���*���3����7��.h��}��)�n��]��-W���-g��g����ߑ����l�� "3��w��t�\?�i
�ȁ҇�5�c\�T�\HU�v�����Fx(Qw��zc���;!��j��2�Òl��{s���&^j�S���LB���z��U�jKo`)x>+}%���烹�<m�3�Á`O6��O��w� Z���~{f��>��i�&@�y˩�		�������-�f,�"H�vi����HN΋��h�E��(罒<ςߐS]�-��	�Ǖj�v� r�����P�z�:�7ҷ���	��Q�ϐ�E�hu�$���@�c�t^e���ީ᯼����?G�~�`��p!]� &F�Df��ey��R$+GE�Sd�9>�� <�pP[q�v��oy�r��iv;t2�ꈠ� ��}�����$���k��^#�׆H!�x�:Z�7؋\P��v�Rez|qT�}NdS��C���f����OG���2 ��ܳ޳aZ���u	�U�%/%�X�;�;�3e���:����dM�ʾ#�9���|���\�4�����P0���m���������w��"��t���q�^��2�b���{������[��:&u]�犥*���kI��f�wU^���	�ʆc�n��P0G�U����g��x�nd,��]���$��h�q^�_3ށ9�N}�#
[
����^��}h$zó,�6�y��s�ʰ��|�3>���~�y�P���f��z�/$�����_u���F�)EJc(�chw����FQ�Y}��(A�d�	�ڽ��Q��~�
L�t��3���J y�U�xS��Rg�t��?y	�3!֪;q�gWr7E�F��� /ߕDVo��g|��EW��@0f-���ȇ%��K�����!�Uo䘗7�Y�Y��]d0o�v؞�G�Bm��5�<�8z��䶾j���hp�0@]v#�5[vC���	�:��PQ6��yN�CR'K���6�%P�����#�m�.���=\�m0�_�j�Z�� ���3
�4vbq����\����e��g��w��R�v�>
�J?X?��o^����{���&c�6&% ��+WY���Ȕ��qX[k"�ȕ��AW��xƽ�����G�� �&�?�<|��?���`U�_�[�,'��צDk�bֶ�*�|��1��2#b ~M)Br����OՏ����{O�Q�0:�~�$���:��Y�읝�L���'�U}LIs���kGdd���zHk����2�PTjàհ��,�s8+ת�AԮ��ճ������p�\Ѝ|nzq�W|��؊�;�Z�ak��7��� 0%=���#�G��! *�5��	?��#S������M|����*q������;t��ʚ�T���R�~�Z�Z�)A������k}�f�|��Ddv�׿�<Q�	��S��f�<,�|�s��x[�*Br9���+g%��_��c)�`���}��%Y�@QL��>�G���	�}7+�~�i��2֞:Q�*,��k�e���7�s�TEB�s�K�x�H5�1П��##>Xѻ:k}FLkG�IvM�y������{~�>8�i��[��)�q0]��[�pr�>uQ?�D�O�>:��^����?@���A?���\��ᵭ��ţ�u<��^? h'�'Cg�\dɦ$�ݩ��i[�%� ���Ĺ~�s.�~"��/ZPq�f�>R^rT��q�/��b{����k	F��|c�:d�C��1�����=J���0m�d�\fUF'S��7=��\=}��������`�/wxN^@��ݹ�`�V7,������g���s
V��2��� dh,i\�c"k�s \gK�Ը&6�*۵i�8fLQ|F螫�Ȥ�
ʲ�qc���p`!5fՁ������Q2gƩ�s��J� �^֯�=����ƆI��Ugj�����Ï�>vRT�}���u���,�	7>��,���p�p-)k-�sY}�~m�1���T�ο��gcQ�Rh���"�S��DY�U?�i��4d<L�����2~D�L��!�Mܔ�G�S������n�Tﴘ�By2�f9�1��N}$娩%�1��=��膱6 �*A/�9�ۭq�P����B}�R8�Ms��'{�ރ����M��,�F��C'���޵����u8X�-�8�LD�>�P���/�Ĩr���")�*�+�AF�V~�@V��Ȭ�\��lÎ�{do�Ƈz9Ӷ���4k^�k�e��3]t�FLӪ��j�K��?��۾�v]?�_!�����A��겨��mI K.���u��F�QIBS�Fa(���C�A�P���Un�s�[�W����k	��f�k���Z����#Ԍ�;'�?V/X0ď��̳�bz*kC��"���;�W�o��O1B?fQ�:f���G�X/�`r}I��ڋP�* ����.���y��!�~�dfʞ��Ta�9��������oqx_Rc�ca5���i*���Kx�.Z�L��ݭsa���y��FC3��8|�Q�ŵ�hO6�%�I��q��c9��$�P�����!wCd��fcx`��p��o6����}�}��>B��:IJ<���#��a�N'�v�?�04�i� �5���
�jâ(��9��7s����>��\����gF�T�����)B2�Ө�o����\6u)E1��b"�>3JG/��#;���Jzމw7x9�MU&�2ʟj�+m]6%���c�igDzR���Vh���.3g�>I�a��
%�jxɪ��%V:�UO�N(k����X9��V�^ ����~4�o?g��g�zdAk=�p�D��	�j��Ͱ�X�੫�_I�m��C]A�ƃiy��e����$#"�峄U_dmZ�H����S��V�=�����0��߼�{ʘ���K�a�FB��*�!x���g	^@6%��)�`�����u씳�r �-�9��-�[����:�v����Q&�?�M<�|�x�~0����=*�Y����2�+u3t��d���4��m�ٹx�H^�_�s���.�krG�7�%�`-ϑ{|��a.��ݪ �ULGf̵��\���H�!6X��,Tw��_�G�AO�D��"v�Ό(ޝ�?�28�Zy���6+2�W]2���"�S.�0��s^���s�/o�<=�����8�
�L�J�q��q&���sn��~6�D���O��҇���4#12Vd�/KOWnwǁ�@��O{:FLX�8j.7�%��L(�%x�ù�p���>+|���@�vI�|F�XKKn��`<m/���i��Tp=1k�X��vȍ������M��GL�Qk9��!�.�\�\J�蔵z�]�=���!7�>�f����n�;����O۝�.7��!т���ԏ�����n�����s�}�e�܃�u�����ޠ������=�jV�k��ڹRZqs`N]M�P~ì���d���,>�P�?Qװ�IΑH�Y��*��Q�u�� �;�
y����r��b�f�n� E���tt�ІOռ�=���>�Ĭ�[Y]� OQ��ax�Nd�P��yշk��3������+E��y/�}+#�{��餀�V)�5��}�s�T(Sv�Jvaԍrc�d�N$��{�� �am��Q��L�pc^$F��ť�x�T,g������ک(� 2P"��X����+�ǫ��Ե.��Yonb����E����/�B�\��}�,���#�L�py)�h�Aq�r�u���"CaW�' ,���\�Pؚ�>����N=��J���q�B�����<�ή���x�G%}m6JkF{��N�r@�(����$��^�%@Skc�̓���b��=�</�yP��R~+,)�g�M�!;?�i��K/;�/����.��aD7�[�Ѿ�65�("�fU�z$���K�1����)��lsZ�7J�ޜ��;�E���q����LRnxOP*l�R7�.��>c�sJf!����L�δ���
{����ld <�����T�~),C�.�fάρ�8�+/Q�������]��-� ���?�D�����(E�5dU��X{��+L��#�	Ґ�r�Ig��{b|���s� k�!'Dt~�@����L�ue���݃OJ�ډl{�KPo���Z��~WkL���g���.\����S��A��7��Wش���D('Ae�YG�����g8T�S$;;��^���/,/c�V���m�~r}v#����?��n��H�(A�ݬ=��C���0�>��*J�߼D���3����>Jla��hTf�!|�/����-��1�sc�=���X�F�3"��ܶ����;x$�g�n�����xW�!�����&rx Nw��SX}l!Z��r�J�7Ld9��vh�͡�.�7�ɩ1d�k����]��P���*S�o?O�3t�䱎X�X:=ɑ�	.r�n��@W�UW�b?)�^Y�;I���j�a}:F���م���|}���/����~�y�C���;$�%/�����.^��QQ�.�G��2����M�υfy�4���!�}>W��kz�L��	�vn�Xa�~CP]*��ύ*&�Va��׾5�HR#�р�G�#��<!� �dT;PG��2hW���y��@55e��ݦ#O�{��`�@)`L\3�_[��B�;���	�b�O4�Ƙ2s����1�r�����Cƽ1� @���u��pI��F�ۄ_�ǨU�+z���{�U�����,]eѐ�I.�H��Ph�VR޲X*"��.�K�e�!f�[��Y�="�pGSCL��wrv�u@�P�Wc��P(x6�:�Z�sM�j~!˘�KE4�/NB�;�Gi�y4�V�� L�Ƈ:��4�8k���k�u��"�Ӧi`���Ιꅏ�h2�j#:��h�p�R���UO�:��#K�9�v���yN��:�����Ν������.�Oni�ju�zG͝�D�2�;�6g�,��q�uj,C�s�32���)�^bp^N�t%�!�#T!���T$�Vt�k+/�J2`���P�0��-IX�#z��KpY4�2Q�+C"����Y��q}��k������+˃'���b��4Y��4��	86�l�߭!������  @ IDAT�ui��h:��9�L�h��ڐ>�����p��)	�i�Ql�Qٸ:�)�����2��1-)������{֜X�*��؂$x��� 򚢎��m�F<���鉬�C<%��d�gk皡���@Sã��
�
�v��?Nƒ|���,3(��ޞ_�b�8Ň6�)�dƹ��@�]��\����Aߨ])�Z/b����9}~3��d9ZK�:��`���&�W�jo���*���*�W�����ح��$2��и���V�:Su9 mד΄=2D^�+Ļ=�'	�_����\�o�Y�<X'���񇒔	C�%_n<�ujO�Y�k������w���B*$�ad1$+�;�=  j��1(�r���[�zB4$>�l�Ÿ���K�0h6�:�忔lG˅�B􈀡����7ah�"T1�0��~91���g�#,���B�)؅~�
@�w�=P���zҫ���W��x����!J��Sc��S�s]�2��z�~�(��0L�ѶDdOЀa��"�)��FF�i���@ߴ~h]1Mt	[�P��a�Zb0�W։,}v1�gAZ�E��@��G�F?B�;e��|�� ���E|�ޔ/���	��Oo%�S��jgNDC
N���z���0"������?�|�N�
4ҵM^�ߦk�칶�����,d�G�S�*WпA�i=����J�����".	��Ca���[n��`�j��?���Z{3x�� �M�t�h���Ƈ����Y7j�zl�i���Ð����}v�em趾2�a�������.]����
}�p�7@}��N�[���OV?�V���5�P��>�w����E(F��x�g��,`��c$0w?�>VYOB�	�qq��lL �h!O�1]�~?Gv"��S�L�vSҵ�5QHG���qY�1�pOU�?ܭ���3��+���E�;��A��x���n�3~ګ�]��:���p@��@�p��$i�5�Wb�ÇkS�#���K��_�Ux�k��� Ff�K��7V݉ (�����!��7�9�V�3�̔ߛ؂��?F ��1�6U,)W�c�l�$�bDp-�܉5k6�krU�"�\�KT��:r���|��N�iJ�ڋ�+�$z��Q�-N�H��󊆳ʳ��Wp�3���8]7ӓ�sS��N�q��d�rb!:Ip���~��G'���Mt�������'�t���1d�(���\��ns."us7��E}���mo�
�9 eB�D�nk�z]'<�o�A��@X4�dG�H����		��p�
��A(����⩪V`ʝۨ�SN�yg����(V��a=��ZX����/`�D) �PkÌͭ�U$d'�b��J*s��nD����Z��*#���9o0G\B�`�5<(�@���@0{�կ0&���b�� �c�p���~��}(`�	�%�+�K�,?�C!l���4Ã��~�Ǡ��$A�ϨD*nx�)ة��E��{����Z)[�{/I��wNíΈܚ�J��{��%t�{�T��%�_Cw!u�C@!P��u2���?q�����b$���s4�^��HG's��'�_��e����9c�0�9�����0
(+�=���ć��仔#N.|#̓��kE��8���)z�| #$�B��7�O���c��A�*���f��8���_��>��n�3s��톍[�TKdȂ(������a��4���r�v����={�mi(3R���~볟齘o�i*�E �Ui�q�1�p�s��0h�5�S�Е��*K�UlLFm��B_���V6�*��Z
�!a�������u��R���5vW^�z� ��R���	�������6����3��Yk������:S��;�ā�ϣS�V@y;��_�J¾�4���i0Q']�� a��	av[���O�	��Q��I9$��������쭩��[�ݎ�)�A��"�n[6�E'�<����q|�=kz�+~�x7S�U�5/�0/<�3����4��x������.��8�÷igX�y\mY��+�@�94����HG��S����>�a���Pk5��,O��W���SW8��aB}�\����\ה��6Ĉ6X{s���Y�o����Z_yè�Ѣ��֦{ZͅW�0C!����;[9�h<�k(,����݁M5:��vK���:��8�$ýk��VK����^^�*��[[#�|b�� ��aNw:d=��-�R�sY��˳<�;�A�.t1�B `����Ի�JGX3bYƇ%a ��6dO;�W���7�ϟ3��=�p%t�;S~v��Aͭ���/�&�۵�����#f3&;�\=x�'L2��[�~��Ѐ7c��k��=��c��	��,1��c�ynNx������j�P\4u���Y0;�u�A�L��{P{�QAT�>���w���d��1�Mpm�����I'\��y'����Qd,(��jKģ'-��\K�!�p�q��X3q���vtF���զ3�`Խ@H�c1�w�t��%E[/��fċ�-(J�gT��.K�;�"c%J���,����cx�\����[����`(�C��>���~'��h|�Ӫ�E��2H�p`�^�8�)	�a~�������R;dp2�c�3dV0�l��=kT]�__9������M���x��q���M��3�Y��A����e���rcNoO_�� ܲJ��\��r$� ���S��-��ޭA�����W�xq�w�X̣ �ޣ֌�z��nQME�-���� Q�
W� `�i{����Ǹ`ܘ���~m��`���7?m�`H��yC����q��B�Eؖ"�ٝ%�����l��T�A��_vz��Dq�"x��^-Qi��r�by��-���P����ƫ�!�F�x���%�'
:
{�;�J�y�k��w��$##�չ��E$M���*׍P���E����"$7�{��{ƀ�����4�8���n�����$Tk#�nMM$�ɮ���~�f�3�~T���x \��B��0x+l�ƻ#�ne�xq������Ж�9�#Y��:�r����pN ���oQ9YO���><[���`}��5z*Ozq�Y+�O&��&ƈs/����ӡ���2=��O�����g��Mb�/ʔm�(=�$�ui;����(���9�`�(�҈���]1�*>u����<;�?�!�u�K�+����5~HW��l߮�R��܆��M#"�-�ʶ�]�jk4V%�YD��X84%V��x�?�{�&G��q�V��*2)8�O���O��u�W^��f�ň̋ϓk����aI�$K��D�C�@��� ����ط�N2i	JC�F�p$d�~{8��1��c�ݓ��g�T�i�!P�6����ȰL��V$�O��g\�uVn���F���p$=�k��E�^��h(ŏw�@���p9I��v�Hp'�=w��й^6��ME*GN��}64��k��f�D�3���04�|,�Q#/�n�O�V�tu���B�O�n+~�<����h���wE���o���qS���۹�f���'�i]��������{����!gS��C���fϖ;�M\���q�8�,Jϳk�Gf�_�@	s7=�2"�Y/P�0��DȲ��)��N�c?��0Xz[���S�5���$���(�R������"W~�zZ�tx���0��~�����S����q6�����.HnAI��g\�d�������p6a������1*K�:T�nm��<�P�i�f�`�s���"Q(!��/�-�:m����3Q
�.OS]����O�uS�|5�!���C!G=xv����0�~�2f�p�gFm4��%Cx�e��:�ŪB3�	�]�\��SF�	������� ��W}ǣ�G�cxFc�@��Z�>TG��\)F�yb�Έ��"�x4��%��ް� �rJ��A��/ʃ��VW�.�q.}A���5'���,S}���ǅ_d�Z��ǉ6�<���Q�Iy�U���\���[�~�&ZU�� �)�o�qe@�i@���(�tr�J����}CĆBX������Db�c���(� 4��\���'�#_ai.F|�Y��3h�? S�!0��V�ic��q/\�1�_;�s�p�%�u�M����������1$ƻ��z�ѻ*��k����5b�=j��;-T%|�6V}�0��+�ZlS�R�VP�B@�%�o��0 �?����6�y��1{kd4�+�����0Ƥ�K�aq+���E�2��J��_<J��r�7jF�`���MS���~��+�8Z��p�F8��[���q�K��~�i��a ���Je��$�]ۇP�nD�����nXt��깾���۰vs���6V.���Q�݅�[GR�g�ȋx�6�
��gԬ�	ܞQ�Z.��7���38`�q�s�9����yko2�Әrp��S1��x�`���n$�'b�E�螁�|�}5�!m�z�̓q0��{_�p;���j�^�6!�����������1�K旘�����0=}����v*�W5.hgE�G����H��{E����b�a:��J�1��+b�rۺ|-ӟļ~�PU��g����%��f�&z�݄��"��9���D<�>o�p][��!j"�.����0[?��H+"�#dd����-��g���c��~F�W��O-S�#a��v�ya���hv`Td���&�9�	��l��D���7w�<�l��@.��[�R'Q��G0-O�B���� �Y�� �
�6�as��SH�fT�w'Żq*/Ѓ�wp�2ʣ-u�Zzx�Q�fgv�QwР}_0�W���:�l}���g{)���g�P>�㣋2���B��}{��6���s��d�LF��$sh���`�~G2���o&3�5���jh�z[��=h^�ȶ���-���]h�.2��GO�;�G �kt��O���P*��� �a(W��j�����۬�R��"d��Vo����������A�tx:�	�~)$(���ۯ�G���}?<�:3ƨ�xS4��G���&��WK�RF a�.A�<*o�p�x,^�'��TH����1�qXD4e�"\FG��#1�%!���f�p?�զ~	km7:��^��	��q�~`���T[�(���Yx��{pH�/�$?GA�%��w����4H���τ`�����?�OK}�gheG��*��{�]a��Ɋ���W���^�kkQ	^F�����m�;������]F��
�d��K^7�&��2TQ/|	v ������W��a�����K,��m��0Tg���#���l,'��P�\�xI��~�98U%#���a۔�V�:2�[�@�O+��W�nIR�ڛ�}���c9���{n�ϒ�W�Q�k	`�tm��$���� vg�'���ޠ�>8ߝIIQ����~��n�����aL���Ĭ<�� zu�KV���3�f�8�	B��l0W��T�$���F�J��H�p'E�@�$�{�X�ku�O��n����e�se6E�G�+��bO�h�FV��q��ʙj$,}�C  `C�Z�X���\��)XC��Iw}1V����Z�x��aK�Or=j͵�ڕ�06���[c�K����`JJ�Z��,B
F3I�FhP��5�'��V��:�z��-���ӣ`9�U�2k2,����_�c���Y?ۖͳ{Fr���f���uq�
`���o
}�%e��mO�aV���N�� �G���.���u�m��*z���g��0'og�D����k�`�i]�@�?�K�u�X_��������ۋ*TKٝ,�^��L����bp�!y�gy��:����!���k�F�V�h�>`�ĸ
��p@�*��̷.���gb�0��`�S��fÃ c�f!I}"�Bk,�y�����}#B��쮿����|�p+E�y���[��ޖW���pr ��Kq�n'T��c`l}�N���G��k`��P8�L_j
��C����{4"��)�{�k�$.�!8�u�����16��v�K񴏼_2�D +<�y�Ď�ߢ�p��ɇ)S�$<��9�nxĦ�\�<K�g|'0�����ؓ����6٥4���=ѡ�_��j��J�[ד���r������S��K{{�5ẟ�be2�mQ~�~��B��S�� s�[�v���cJֆ��G�x�/3��o���Dv�'����æb���[f8�>���3��[T��9گ��23�w���딩zyؔ�y��'��<�K �G&m�%�n�5tsI��ư�C�Xy��DwZ��� �-��#�{P�Dk�c�'�^��-��ѯW���`�ל�s@��T
���k�NNi�P�HxdL��ݝU��+��vy��Ix�3�@T�H�g�þ�ڇ���꫿漷&���)�V"�����kW��i���bos�6���W�wA����|0axu�	� �>��}���]u��C\4�/?[��N�k�.�����Dr�>|)5cqr @;���^
�J=��1] ���I=�&�O� �ѻz� �є��<RS����ȼ��=ېb�9"�>�P�m�!��P�#Z@V����n���7�9��Y�@ �
�E�3p������K�Ur��Q�'��B�������"��.�P
�3�����[�]�{	{^ymT���\hb��Z!/h��9Z
�xñD,�����;��͵�O��Z:������܄�ϫDj�������EDEEhF���q�l�0'�A������D{ֈ���{d �]��~I:OB�eNͰ�����N���οx嵨E~8'C��	^Ӵh�5@�6��e����DH����x(p��3�2A�y<?�^��nƐ[�����q
��>��_� �X��?D��%�j�����iOJ��`S�G�8`�'�����Ӟe�#�kSF�ԯk4p�V�LЬw���B�y���[WE��ZڠF�0o�l���O�y�� �U��Ԅ���/\�1R3��t��p<Q��Q8
��8]G!k;�E?²��OKn�bxWm���9���A*����ĿBڬ_x�]	Xw��H����͹�7�rBw�2WA$?�r��(l]�M'���s����oS�`�� �?�@~�a:<n�c�K �d�d��п)3�5A���ɉ�,�~��8��E�~�U�V�r��	�73�1���ɶ�5ZXɜ;(���<d_.�.��� Y���o�r�[�Hp�1	[��'������R��0jVn;����U�ʔ��!��b<;QJ���1���p���}6k�ڀ�(<.s@S��݄q�>� _3u���� Hx��>3\�8E־D!&Dqo�Wn�Jե�)�&�� �Zm?o��N2 ��@l)p\�N�	k��|CD��s�un�h5B��Vs6�g�B$�I0΅��u �R�3��_F��$���_P,���M�q��ϷZ�L�nfK�۷�6&c�1�htm��co�we�����g`6�ݝ=�	8g�o��.j������@ʡ�v~nkq�a�i�M��ކ�q�h���i�ɢ��Z6���h�;�8t�.ņ]��rv���S�c��y0`F4��UW�x�s[���"���U��)�5��]��%�K�Ç䅡?C4r�[*�	1`fi\WG?���Pn��t����o�=3d�)�ͺ��Bf��DW�TS���x��˞�B6]���{�ߌL�G���8�視eF���0r.0����!,�E�P����1�λ�᯶���p��*o���hJ0�H݋(�mL�GG�����!���6VBe�xJ���ϛ ��8C����N�=���[����c}��П���}�i3W�C	y��G���uYO�=�/���Q6Ə��+�&YDA1l�^97�E��xB���y�t~�F�..�,Q9%�1*�3��A���Q������6�u���|�댮��9^�V�_# ���B'�X͌����+��$�h�����C���OH��q?x���R[�  <�B[Kȷ��h4�����-+�f�&g�jS�FF��f��~ O�;�0ȷ�qP��wR��)�U�Dp7�U�.4��2Q	�z
���g����GS��))52�
o������Z�,?ڈ΅6t���6ɒvg��;|����b��n�)��_�p�~�VD�7�U�"�vU��x~�p�9�dC��	�������f 8�"�����:�vAL�#�g>����y1cn��C=���������3L��%�c1�u���~��o���͞A��f%���u>ck�j˥=��	���Xm��O;�_8W�Hԯ�ԓ�U���;4�=a��� ���'�!d�ˈ��qP�%.km�S^ �e�fM��TM�9ۙ/x�`��)?�tc�pưY;}A�Ѝ���J#
_�G��c4�3v_v�`l�o�ov���x�p��R�)@u�E�·��wy�vm.�6ױ��YSa�!���@Ft˹+s��`�(�xLa�ط1����o���` c��ʌ�\C~}jkg$�>���)�(Ё��#mwD@���i��)4�,�LZn���oD$d��j�.��Wy���o��YG���l7�-�W�$E!�"�ma�o��O����!�rSji7�w�M�6�B�W�n�L�S����%��d(����I���G.j�>ͥ�c�tx�o"��>��˫o��um�`�w��06 ��Y\�<F�Q=�f��OMb�a�~|!F%Pc6�Z9�a<#��1>K�s�b�B�xre���㑶��Y��-gGb�"FH��pl
�����a�傋���Ո�E)
;��h�:�?o��/���3 ѧ�rÝZ ������c�F�PR�C�?_����]	.3J-���b'5��a}�~�= @�D�k|�"�G�L�*P�<�� �eY���J��^��b2R䂮=��h��/F�(r3���^��7�-	3�$Iy���>�N'l-������7����锬���s��j�:�#��d"��X�t�\��W�1�lw*�F_��y2 ��'V���e�_�yu4T����0��f꘱e����;�>��ѫ+~}���S���2q3`v��D�sJ�M�w!%
���z���"1E�:����ݭ;�܇�h�����o�ָ&���� �q{֞2kY�u�����u��QS��m�B��9�hB�Oe6V��61f�!�WG8�+
E���-��"YÙ�)C��7�������"┼:��%�1��H�iSH��9o=�U�7^p���0(����-�N����=c ��{�c��������w�?�j���"�o�@#c�Oʜ˝���Qm�K��Q�hH�f���k�Fߠ}��#���#l�
�	e	`BD�n�3Ve6�A�Bk|�Z�Jzk���+�΃�<\�'
�9�d|��zl;��Gٺ_�"�� :�s����v=�G����"6���lShImp^%����s���r�!�Ɉ��㱡M�:��3Q�9��0�g�4ɂ���ź �)v�i3Q܌5`�����p�caD�ȵ�8>�}�H�G/��G�(H���^�`I��� �"�Zz���6�����{�r�3�5%T� ,�z���\^����SB`������5}5hu"&bz,��x�8���e^�)A�I��>#�Pn��F�.O�@l�6z��� ��Tpeø1����
��F5=`�7��ch�6���"������F8-�6��+�p������������_Ő�E��<ƽ7�zxo�M����Lh�h��c��1�7�z��g�/<� hÎ��aVQ�Ӗࢍ�urF�����s�m\�<�1p+S4�j�?�+i�lx���ͧ�볦�RD.ќ ���9;�||_k��I|� ��+/�� F�yr[�_P�h�Je3�7Qe�l�}���l<����m�Noؗ�9{r�a҆�q���mfB�1>���E���p�"2��9+�^}�� �R�9��]����OUo�[�E6A�a>��;�RBm�m�]�w�It�/Tn2Ώ8"�M�D�0��j���S2M4�7zT6��!\���C5�/r���@�'��ֽ�������K�;'��x^�G������?x7�J��i�k	�:��nS&/00�,���|E��I9M��.beM-���ϛ�-��ӸW�d���'���	�����}�3OR�-}$��p���[��)���J����،Q������nF�ND��HH�I�	�����")�6o�����EB�7�XtTS1Ӹ8�N�g[�}&�Y��ֲl�^���ʿ-v��ϮՋ������Q`,�e��2�Ţ�-H�b����?��{Vi���w���`�$pDk��d@]��"�)�h�����E��
�z�ZE3�5��>vh�%��:R�0�w�����z3��L��"��5>��W�⬃��R��o�A�u��C���_�r{���&�=;2�o�� [��}��F+��9C��wZ���\�wZ���
&g�5L�3�G��Vтa����%�F���g w��K���#�z�E��[��\.���3�@�ڹ��h��Y��X��y�z����a�A>��\b��H_�{�S��̾�dw��Ғ@����!��=��?�C��+��/����qS�X8�d(��$LĬ���x�� ���!0F0y�<����P��W4��y
ys�J���PCQ�ּh�r��aLG�(u���b�B�`!p�����u���eY~�#3"2r��v�6ƍl�%�B<G~�o�B�,�hh��CuW�C&��o��v���s��{�5��C����Ǚ��A½`�lCy��H)���d5�/j5)M?�[K/�6�.�*0�n냒�|�H#u\_{ *�������H�]A��gk����'un�,�X�߈.��i�<����]��5�D�[��$���c�TL����Ȁ�>u݆�j1"ݜ�S:�Lm�_�0�������-Z$�fGl]�}<3�E���0U>�ad,��+�.1q�.���<`m��Q�O�7��\�Q�x%z4��ދ���*��ᘓ�>f'kD���o�E_k���c���!9dd����n�i�N������o��BѐI8�~��G�d�>
���C�1u�S�t��9���K.�-v/��gf��1F��7��if)�p����aQ��w
�P���88x�-ֿΐ0���g� ���
�9?ϋ6Tk�u����8��}3
��
wk�9�|QVv_��y��ytt
�?��O;/���"�(@�D��wp������O��=�v��w���*F��4�F�2��E�[W	߯w?/�bR���3�^���ސt��B�.��P9����Q?��W_�p�t�`����]S���t<OF;!�m�u�Z��7��h+8c�|r�\�+���e�	G�лd0�� �x����n�!�o�ޛ�
㛣�8��Xl��TzW=%p70���H�}C{|a��e���WY��[���Ww�*���$��[��z8p�S�7#ap�$�ғ5[�D4ϫ���Y��/�����c�!�W�VtN�%�*��~�`[r�����f�В��_� ?�
1�`�e�{Bܯǟ��P컿���(�t�(�=�!���^�£����ө�<�;7�����1J��Hz:&ɝ����� ���1�S�f�:ܐS����+��9���+'���Z���	K7��F��Vb�L��QWqV<���<a��녳��Ř�h9������'��10L�v�%��1:.|f��uO��ʑG���{)�imu��L4��|����΄�����ܟW����Qtc)�,E����Lng\�s\(o����[�}ח�������C��/����4]9�g�a8�Z6R=4f��k��\X����K�M$oV,�ѵ�n���T"jqoj��4�1�tQ�7���v�����c��烖�-���`�l8\��Ɗ������m��F�GI�vk�� rllm��i��mkL4����D9���j6�3����A��f�X�嗿z���������b3]BB3��H뙒�P��z�v��@F�Ҥ��3�	�^7a�Ĕy�������(nƠ[���#ݵ�-�]�c����s����)�u?V/ܫ#���Gh��"H�	Qh��cY+��;ܔ"�O$�����ÁMᐲ�y*�����҈$�2Z4&��;��A����������ϗ�e�1XZr���Cv��g�u��5�T��R�GD������(��V�1�MC�T&g�d�c�A�7�pDL���P-�S�����iß󡸟��:��~|�e���t$�����e
.���MkO���"�"�#�B���c
ѡe�߿>�r�L�j�+)ߢ�/Z(xc���u���HUN��C���']����{���BH��S��2�%�A:�U��m}
t߲�������ۦ�x��bNS�����X��&jEU��'�m�3N�?ENFŵ�S����o�x}\G^�/����y0��u�QR�	c/Z� ���ʋ�G��p��%�[ˌELDz�a�;cH ԑHˡ1�9H��׶b���Q��Ì�D�c��O1�&(���E�ZҾ�^�8l)K�1���C�V���?�cf��\AK��'+��x�I4�4\�dǢ�FF!vNT�@хL�<Uq�㔦<i+�Y���(�^���4�qG���N�?���ZX7���@���#�@�����d���%�@hXD��DY"���Se�˫����z+����](��A���\}6d�l_E;�H���4�,z��1y���?(�3ʘ��������0��(��M����x���w����f|}��w��t�.Lό�ГK"z@o�qR��j��s�f9���-2�;��OE�]�c{,��D��W��۩h:\�ѿ��=��7Y�,��+��f7�vSQG^��BS;����/~�rk�ߔ_u.AV�ЀLN	^��1/��J
��P
�ew?c�Rq���`ۦ��Kmz�)�c�#l٫��31�o�m����C-���˯�2�P`���l��mKd�t��h�fR�ʑc�z���'þh(��fJ6\���S��l��������B�E)sU�OX���������?���jF�
����:DDp`$���zϠ�9����Z����nsVx�/Jd��`�g��0�N��ʼ�̇��KW����^+���fȀ2��dhol���19:�I�mE�_�	��W�̈���^p�^�s����Q��� ���4x�����t嬫_4'ڵD~����1�x�A�{�ݞ���F��A����W���+$FWzA�����i|��9&]�[�gA��+ƈS��\�����h�#��,gj3��Ѡ��U��"� �8��3���1����)_c<�O/�������{�_�w���&c����O��׼�djpS��N���y�k���<����4�+7�A-�p�ɰ�Pm�-�^֫�����C��Z��OH���|x>D����"�K`���R�)���Dw��We�kSC��\�����c��֚aWnI&�FA����_%(�ɨ���*%��oO��ѱ5 )�Z8���c��*h3=%�[WnȠ_�E�S�7'�k�ѥ50F���S�V����ZV�9���?��Ꟗv�V~�1�@i�Ȁ� w3^+A�e��l��>�e��Z��YoI��ϙ�j�	L�-މ���@K�2�;E�Q�����چ"�|��4C�6�Z�Pd����_�u�=TS�9x;��s@G"�.�/��"����sGꇬ��"$|���.��6�q��Н��)�{	Q�'��s
��'�p���r�����5�u�,��a��ZIպO��,4�-̪[�_.4@x��"���^�-\�ݲ�cb(/����Ms�2qX�cmD�5bx[�Ho���((}�f`{O���J�E��փ!�3+E1�<�~�.�3#����S�u���A1 o�Ғ�6f�����y�;I�x;�q��(����S�v�h��^N̶�e���;�1���b3����:�A�����RD�ʟ��-_?���+�9��T�=��ٿi�Z�s(g�{�	b�G��S��U(��ED<�s���#�놑n���xo��4���Cx��.�e������brj7�e�E��!Rt�aǫ���V����u!�����Mu����p+����7g�"��#/�ĥu}�nQc8Y�,ɣ�S/8��W͈Y##�п�Z�E�䑳ͺ�F���{$�o<-�x����]��'}D�;p)
ר�|:Mq��}���2�������p��>$'?J���Y���V�8�L��{{�S�q�­�h����Ȃ�?�uF�j�2R�)�0C
� ��g����q��*{_m�%_�0�VeT"%�(�2�'��b�y��%��4j�g�d
�xz'<�_7i��j�բ��j�rwl���2E�{�F���GZ_�l����][��6�«�PcyR����uy�s$x-�ю�s9������n�>�9��y��N��z��A<�'9W1�?'΃#c�7��o�Nӂ�6q�3��!�ּ���(ـu�
@�߫�%������c0�V�<��k��q���9�j��K��\]+Ϙ���S8%�dg�����v�v�r�^��N�_�;�V!NObդ@��0��3��I�Q��l0���<;�S�M]����h/�G��B�O@�=0�6T���-ŤOkX��8G�p�6�^"�>�l���\}��^U�Eq~�DG<�jD�"(�$s&a�GP���Mn�q�?��j�O���o^������/�'�&UZ��$���@^AK����%� �`���7�0Za�E*Z�0�~���L��@(�,gE��l���P�@��b��6C	?8�L;�h�W$���%a{>d)���`o.�J�:���U=Y/_��}R�:F���h�pyv?�-�![(Zx�}
�X�/T5g��W�#$����nIvY�~Z��3�t ���㏷ �破i�y����Vw��t����Z֮U����Hs�0�����C��؇f#,2�\�F��9�pH�������E��즋M�~����FFS������3�"�`����9WO1�r7��~��T��Ck+^v��N^�N7$��FW7=㜴�t�>��9C��U]N���$�\}��Zӵo��i)�����n��^;*�yZ>���8l�� p�a[I���]�p����hK'd��Э�t6ܟi��Ǘ2�/[�s5����A�l/���"���e�����?������?�/�ƼC$`S�4f��d��qO�°�I� a�#�n9�'��Z����8ϴ�2\�J�?�~w8����G��P,�I��n�|8����"<t��C@BB�;�㘏�[Dշ��5:<��O�{;Dd}F]��LA�JTP����#d�2H�R�C)��#���o&�������s:��Wv���Y[�j�����G0��o�K��b��=��쎕����-
�c3�{����b�܊�K׽��6 ����zק�x_�2��_4�!̱4zO'��k��G�L5p{���%��ǿ��N8ϥD�wu{���Kg�c�
���~�0�g@�|g�Q�o��\�%�5�0�	�����pR���+BT\Z�)9�nИ���5��WW+5T��Ӊ���Yg�e�Gp��>�E�"c�D @���_��9�����(������b/V�ա���M1�A&�d��ٷt�D����YC|�p��z���E�0]J6�ԴL#Ē��#�|����H��)ʼv��2�c�����^(�o�Lσ�E��7Nbf\Ԛ��a���XC��ݥy!~E�%(��p�������ak���)���?Z��I謂�����9]�u�!-����xi��dp�č�G좯�f��_6��S�4��M���Ҽh�j��)gC͓�C��r�23~-�\��:��u�?���
� )�p2(ܢ��<�Z��x��c��O*�.��`�8ڍ�p��~\X����P� �AO<=��t�'�VK]Ξx&у ������L��qx�ݝo�v�e�:y�w�Fj<T3:�'���m��<y���GY�����#[�?�tM  @ IDAT��x��A_N��9ޫ�B7�m�,e#[�,���#�d�fF��3�/"�����U�ÙXr�곊r�fCh���HOv>�����c����P�Or�5�������HeœO(�i&�	��/�z����2�	$	��oS��/��6]�Z��c�U�RP�@�۔B�Rd���pz�ZH�PS���7��!��-�{^�2ƼX��~�S�G�`y�B���p���08<
�!��J�=B~�,�+{^%+M����Za6o)_�5u-@K=���gD����ù/&)M� i�_܇��h����y
-�6�p0;�iU�ڼ~�U�7YWZQ�������K�MC,�z�j� ��s�O%)=Ã��I�y+�Gg�����O2Y�%��������˗�E.��mh�ӫ�ױ��oh;I�j����C_���a�k�ѱn�^�`�3�F<Əڽ� �6���b���$[�
��6-�6L��?:R.�O�����VkARu�E'�hq��Nk�I��	�p�ǎ&��F�ݘT��X,
�������ǲ52]���}WG>�S�K���3>�b��~�*��/��ߴ^�w4�� ����a�20	="s�'F���4���p����Lz"$7��O����(�?��W�	��Pt��(���>'"L�yYD[�m��R?B��_�sJ=��N	�@�5��@
��ݵz�|�W��U��3��u!��R����E��%J��<�x�)�rR��,��~7�k�]�-�=O��M^�~[��%�&#�r4\�~�aF�a$0�D>w�Z�M���)&7�9mZ~��Ս�U]Hk��=f��Y=d1%��'-h:|����0��*��?�1���4��3�Ӏ8�AN��W����'Ơ0 j>�ϭ�	FE��*Ҧ%���;����g9��#C������h/籮B��x���P��0��rj�����a�6�nN�u4�}�hÀ&+�)܀�^�\������3����7�?�st�-Ջ7�_�����B'�|L9�!<*�{��B��h0�|���+}�����7/����v������Ӧ�*j��u�������¼k=�/���TSfH�SB�/k������1�!6�B���0/r�$��>�Ю`��l5%��KU=�a�����_$�π~�I1S��X�֦Ž����������<[��Mo%�+]<���ƃ��%��QZ8������0T��9��=|����۠�T���d��N��7`f&��@��r�3l�<~��6�^wNt7j-�4���x�r�|aٞ����+����!��!��?J�T�.�d*�2�!�t�]����Yʼ�E��(ޥƁ���
w/�R�wѴ��Zү��|��4][ɭ�xu��r�X�lL�8@$�{���:��;�B+k^� .<�6��I]�'�q�����fa쨕�l��C/}z�ٚ/��^�o���.�ʲ9��=��MT�7�?	s4��in���d)gP�Rw�us��s��sG���{g�g�p4��x��8�����X]�o��v�1��!��P����f��=�������j�d}� 3��y%Rh�>Q��*
���Ḧ��v]S|Zqe�;���+�V�g� ҜG��O�9�1�fJ�;����`�.��L)��E�4+��<�g�P�v[�
�:��O�%���� �����7j��O�z��9H�ql8¿�����-r�Ӕ;:�%�_4 ����\"P�Q����(�ºo�:�Y�to�qL�i�ߤ_��$�i�� ���"�)g�a�x�L��z��K���4GV��k��h�јc0�gy�;�9�s}�v�]`��>�&������b��Fr����ԝ�!)�v�0}F"�[^��'�Vw�����㬭�|Ct4�	h8�A�f�s��R�r���\>  ��t�6�='\M���!�QL?:%����t'5a��m�.*��c�L���"�Q��$����U�������������W1f�z>z�,O�[���c�e҂��6������rB1}���D������JD-��s����:x]���>E��s�r�{(˓�e*��ΐ����� �����������f�縦Т�4�-�)��5 %tQ�4�us�E�����Mi��#dqqj܄��R��?��L���:Յ�)�ъ&Jwr���24�E0{v�9�Zō��,dEA6 ����P<��>�?S������G��I��ڽ�v�<�t'ET>�� ������ɰ!l���ñ\អ���3���1�������c+1'���T�����9P�������V���'���Jp�?j S�(��\����һOt�3cS�I��A����:��<�� 8��s���8��R2���~�����.Yxf��J��[�mz��ǜ�.X4s.S�dc�覼�_��L:O�jV>�S�) ��� ���t�b�s1���������}��r��r�U73�C���A�@����u�+�g�1�ܣ%�|e���)��ё����k�_�e�i �6��*�7ϙ�����"��o��	ʂ�)%L?�FÒ�(�|�md�9��Ĕ�wm��W�Kp�2n�lBi, !��MV�3�h5���)X� :��ݞV[�����1s������OKh\��Q���萹�l��@�3B��gb4x}+np9�2p@O^+���2�߷@
�Us�[�W}X�t9��t_�U���n�W�!����ȑm0�����7�G��Φ�C�����.xs��ހ����d:��HV��_����'uo׽���!G9�/�[w�(�)嬀e�"Z�L�϶�cz��R��y��W-�j�Ë�g�}��gJf^و�t��1��_}��k���%��鮇2���؟�!s<S��J�O!zލ)�@`hf�pB��7(#��BR=>@���YQU��	w�R�\�lp��0F2Y��B�Zx���1�'�~ǅ��0����|��]���z9Z�����W��p(�k]�+��%�Dk���,��'u�����E=������w0�tݔR}��L��~�F�d��l�S���z����Ӄ�������
&������\m�����P���,�+3#I�^;�����9�d�[�oDu���h�Eed��9Pz^u'�sy]���=z�П]w�q��#��9%�79з�7p��W T�{���ϡ�]�ɷ�:�N�]4��vu6H<1pdH��`&~]^�J�V&RZ���zɑ���`\�ė��g��&.K�gtEb}�hY��Z�W2�Ϸ�o6��՘
i�
��7��7��!jd[(9b*��㖯�3������f�F�
s�]Uݫ��.��qx��	W;�P���{�ǈ���T�[�L����1�J˽s�r�`-q �T(1Ͻcϟ�����}e�KQ(
p�_=�9 ^^Co�C���z����Ϟ����3úS��>E�ݍU��&��fH��2�.�ޘ8�է����㑁YcF�+p@����J���V���A�"k>l������0=jO��?������0���*_d��vV���C{*"rp���)�O9�Y��4R�܇L�8�Lc�[���/:A�F���� �G���l��ߡ�9�����e[̥���P`pG�p`�a�r�	��e?��`��(����F����C>�C�z�E�ژg���e����Ȣ|���F����_�џ�f �y�ċ�_]q!�!Y�B@0Lu�~ׄ�ge1���i��>�<���d>Ģr�b�v
Lm�^�$Xʞ�0֌w������ˮ�[]|�n$J�qyD��S&���E��崙|�ud���"�-W}0{�g�xP�:����c��6~q�D!-�_���Y�t��F��E_xL��i����/�-�}��5S���e�_vb�E	����x�''K43�Z�0���nQ���\E���[wf-=�����+�6�e$�3hTS��ǧ��+��?���	;�؟�V~��|)~�̧~���t�㯓�����յ k��UG@��D�k:��y�%����,[rW�t6ֆ.��B��o�U��N��a�)b��T�B���4u��jQ���n�G0�t����Q1�%t�]��$�W[w�xz�A	���e"p�N�*$a��ǝړʻ�"�V6ş����;F0}�>�	}b���wXM�{&�Y�k����x�������������	czv�2^�/�Tk��|m��6��׿~�xM��m3�3�C���3>�܄Z�͈��<�B�<����m8�O�u#�ut�Lo}�ȵ�����N�"^�ـ����J���xÑߔ�����ۢ��9)�� L��7�E��x���&�$
`u�z��"/�9�"����/��	agLO8,R���+��飺1�e����bZ��
k#�Q��:<��.R��|���� �r����O৵sV��*Z:a/�Q�ڸR��������hw��<�����	ͷ����wΜnkd�r�}?�Ì.�T�-�F���S�Ƴ�&�mo� |HN��7����������?}����u9.Գ�m�0!������S�%ȭ+@���@1&�L�M�<�0i�MZ�4�� g4�Y!|�Ɓ�<�0�yЭ({�!��rkq!�Hp}��B*c�'�0Ƅ�%�p���Y��p���s�$
�9���_��^ZdNY���6�֍1��r:�ExW�[Cp*5�3�j�C׋�?y��a�c\����h��[���~�YN9���g)eI2��&��u�z�a~W$�eR�삏y/���><�D�M�Z,��g���%B��#i@��-����'?L*�EO7����ƶ���|A䍞��7�ݖ&�yZ�xZ�e|�7�d	�v����ʥ�_V�e��*'g[�Ǖp�MR7G�ZE�|�Z����g>�3VQ������#/v��ץI��N2!�2~����֣�[r�8�d�4&�����}�eŜx�u��C'�-�A�����9�����(@����#Qv:UA��4��W_������߽�)�O�B���|��e�"���9�"5%L��P�����7�?bc��7�KP� ���p��Z'��ct�P	���xhE��O�6 9��1 lw"���(���]���r�g�6���%�L����[�\����;�˦�@t�:e�MK��o@��W4��E���蘓��P�7�׶�ۍ�s�3��Zu���B���r?G�{|]���L�)���:�%|`��+�E�,lvJ�O�����{��e3�(ulƪ���
&�չ���"��ѵ
��kN�l���_����`MB�jα�S<����x�����oG�O�i�=g���p0�h0�s�7n��l+�S��/b��P����x�P>�c�砜�1:�(�;P,k�O��rE�1�9���3���@d��䱈%ֈRԯ	7���������-uz�|�����?���|-��磐+�L�w��!��?j̮r�Tf%>ֿ�X��6ASL幞i0+����_b�A�$Á!dk�W5rOi7&n��)G��%؟8�Q ٝ)p��6�+ڰ	��z�%��+g��t��Cm(����K ���U���P08�РK�·���ѕ/��������.sP�Kyuq��"�V�^���cy���*�Zd.O�;���6���\3�Ep{��H���yq��d�=�T^�S�+d��;�V/�A[�/���l���с�Idrǃ>{�)�o��>��K�ᖂO?Օi���6|��hM�0�wӼ��T�C�9�{/&�<Gr5��c��Z�����#@y�$��f<�gFH�p��>?:�\����p��X�4^O�Kؖ���Cc��}�!�TI��5
��J`:�����63�a��[W:��	;�l���Ng���79ǀ8-�;ۂ�4���,W̪"E-S}<{~1J�I�ys��<Ƙ���^8ݨ�#�⼴jآ�����6]�q�7�6%��S0SJa����"�tGe�1�.-/G`J���(j���2��:y�'!���|���.d��S��f���
8�)��.R�˶qNqǕA��Cw[�Q�M�U!%��""43
6|F�!P��G��;k-��S鹒oE>��G�}�_�8��`�����.!=;'Řɣ�8C.���`�����G@h�[>F�H�E'��Y�u���/���;��f�������������x��f��+R��~��SWԖ���zQ#ϵ�t���*`�f�@pו�8[y���?#8��?�4ݱ3��]��v��Ʀ�׺c`�����|���s�Ĩ������h�U����NOѮ$���l4P��y\������1�������4Z�q2"<�t�DQ��f���P�����]���A�
jAAB50�3�����7>ol�@׿�x\�Q0�'_���7x�7�3n�C����y��jJ�39,�ѝ��x���o�+�Qya�mj�)�.��b�p�,�����3A4�F�D����Gz:J�QM)4����RWS��7�}29�辖VԳ�q`Ա�Y$�S��e�˫֐%��<���]���k)�o�M� �mM��!ʿ����f��m!��7`�Ky�{�E�ǐ�Ϙ蚄w���J�??�)L9L���}��X��pr`�V�	��~%�=��ݜn�
��������=�6��p+�L8X9z'wM�?哞$W��-����`�8r�O~���Þ���#:���`���j���e�{�Ҁ���㇮�{]��f�P$�{sj���~��o���ol����A��v��F@�m|ʋ��a��I�"nkٻ7��#���O�*W`oU#�9>uLFȜI�v�>r��+�[���?$Oh�!�g|]3���Wc&��}|���)a��jL�|�r�c_=�o3ϭx8��)Jh&d�>#im�c8ZC@a�|x*����w�ϺO0��g����=xO�,���S����L)�x@��ފ뿣�g����	��g�(�?�`H_LOZ�}x�{�����)�.�d�֢����Q��gKݗ�������2<���]�ZT�/�=G�a��KrT��FC��s��a�)�C��yL�%�  A�����`1{XR����hb^�AơF�O8�O�G�ҵ�A���m�R��� ��>9��ug=-?c�)wi�����_��1��uq�.��շ�'޳������E������ޤ��������*��Vh�%��:P�Py��<C�{ �,�@Z�k5+�У饗�Lawk�t��B����s��Qxa������7�{YwLW�G�g�ֽ)9�oÏ�r%�-��__�&�݌��k໫۴�X������(�f �6��ԝ�,�î�������0>t/�(O�t-z�����(EV8��#�1�k�\KL���fL`R�tΔZ1pi�W�<!�?̀���EAA�=�u�FNc�V���h:��ڨSܯ������Jh��p��욾����:��v<��X����I,��Z3�Ю�}rX�@ݘ͛pqP�Í^��/�����`�Y�@k���Ҍ��֌Y�ᭋ]}s���<;`�`���x�h��dP��SR��~)���Or��$�u?�����Յ��3^��Ya��2��\��<Z��Pj��`o��P�7�*���^��6�k|���Y�3܋ʾϻ���~�0\x�9�
��� �X�o-�Nߍ���"��)��� ��B��b\��o�NfCpJS������K��Ϙ�h�s ��a�M�"sF`W��cz�e^�����?8�ʔm8r|q`�Q�r}�P�1⒁=�E	v�u?�\�|��|�w6�	�b�0��NC���9��9������#޿mѵe�s�g�τ{����`�]�3�x��!W��'�X�<����a����Z2˱�U�e(kG�¸j�o$�w�Q��/���]��c=%������M�rr|^=�xrb���c�k��c�����	!tS�?/=�o5�C���$y�]K�G�N>p�b8D�����Nೱ.�j�B�N���In�ǼMO��teM��:�z�#j���]���i{����ݒ��Y�O��Ӌ���-l���ǫ��z/JֲnMNMs��H�E/,�'�P~Fq���L�����1�_�Uc0��[�'�����`Q����o!�k��4c�""A%/K�e��%�I�M��Sܼg/�k����"Z��#R��Pk�W��}�'#�=O�A���˸7���:+0�ܜ�V��k�P� ��Sv1kN1������r߷y��BW���w1lܬF��)c(�/�R!�V2q&��#���1LX�8��_tQyi�mL� �7����w-���@u61�j񄷖KT�寜��aݨ�~�i��aS�������4C	|���'qz�o%���lp���{;J�{�X�"���h~����+�u�»Y&2�;z�}c6�t���%ѓ2�/Ӛ�&9��H���5_����k����{����)|��>�z����Hl�۸�y�4MgD�h&?����A�WL>��g9�p�����S��%�q��'Փn��<��6B���/�)�2|�xM����D'5��\#���8T����&y�_R��	�k*r��1����'�p���^9�R#�kJ�f<֎��z�`�Fϔ���@
�(§<WF�=S&�V0�`������X�{2�W�2�E���c9��	��o)y�����Q��Ӑ��&�m���"0p��k�t%���Ȕb��_r��'�k�7�(��m�°|9��=�>��P�w�C��"/t"/'�Gy�Ǭr��4�Zdr��}�p��!�r�H���8�� ��@���gL0L=�_�9΁l����~����m�9�NnG�E�s�o	iϷw͉���$�p�����Z�sݯ�1�m�,u�I3Ec����|�y],c/zc:�A�R%��k���I�S�ka�^�ۙ0J��q���;�*��!~����?�<�U4}y�^7��ݨ���Pr2f��9�n���AGn,�;�e!����P���Ƿј�ѿH���Wg2��gpU����
L?�7}�7��X��+��_��xi���1i]n}��b����S֧��;��� G�_�jp�TOM�!Y�2��9��SiSj�M9�ޜI��P�w�n���|Ʋ�;�6 �"�R�e�"�Y�Z���P	|*��RO1s01`��A�u��*�ȅJ=��U��E�t����� �uJ�	~l�[}H�z�k
��6��L��`D�0�:ȋҺ?C�h��Q-j����h�����}Гr����(B��݀�Z�݇��~O3~�CU��mۅ�����&��Y��u�YÁ�	s��������:�	����.�)cxL�ȶ�OE&t}�h���X?_
�0}�`�M?���U/�����[x�6��F�\�F�W�zF[�SBپ�hP'�����^>��$�Sz�C�B7M\+Z��w�t?۪���E�t׹�9��Т��l�:�m��{b�@�����c����2�Ow�����x����O/~��?�3)�[7 �i<a�0{�\׺D��&�2=BVN�"�HY�s~u}�/�{�b�\��t���R��Ϥ57a_g�/�N[�X����m
�L�d`�C#a�G�¯�e���N9��c�g�i��J��O��n=��{
�U���F��|h�e�.�O?~W8�"���ݔX���/H)��h�E5�IYRƔҙ��_�� ���fy�þ�y�]��3
.!�ӕ����JWy|vfD�{O������%����}�^����q%�Z��@�[�E�dY��y�pZ�q*q��h�����Vn�W���Θ�s-��݀�C���<��;����ӡ�~L�V�������Tl�"<XEΪ����J�� ���B�[�W�]e_���sP�� 7�f,�\��E�݋�Õ}��}�	�YL��01��6�|�����k�aZ,#�=����ּ��X�@��n
�o3��p�1"�cz�$�W�Z\ЦT6���*B,��`�i!i-pp2�2���Q�|Ϻ7�Z��*�i$��aD0R����u��2��Zm����ҡ�3S���^)-�)C�g@�r�qt�i���-݄�V���4��I�ȥ�)�V�h�x���6�F���m��muX�R'�D4���'�=�r�r`+_�!��9;����#��,��a��=��R���[�}c>�+�����?�
�k0���7ys"U]\�+��,J�2���c�u=AW�l�q��L~ۘï������%��ۭ8�v�n֏(&�2F�3=">T6�F��l��c?���G	*Ǒ�uS��Oǥ9��ϽdQ�ё�D����_�u�NG�i��oY�.XkP��������'U���/
��Ɉ�]��*N�ׂ�F�B@�"@Ij+��g0p�~��)��=#���E��S1ؘ�@0 ��2�[i�O�k_�뢜fV�1ݪJy[u��R�F߻��O���/����Z�*�q��|���՜���pԿi4���W�:�X������%�������9�&4̨'�wϞ���S���=Ȩ3���p�s��b��8Gn��qi-���o�.��_�,��8�/L�_�NC(ߣ�UM��_�T�'��q�~���_gxez��`M/���>��2�y��� �˰b�����
o����[# `Y�}˳����+�Њ�4"�h��8�E]��(G�N�����,�&qD���m�q2���q�9��뎮{8�6��I]�Ϛ!�k[�\�F<����"	<�/��ҍ��}y\O/��eWN���r�m�0�� ������Ֆc�R���r�Ǖ
A�
�Iա�iZKG�z#�=�,�1oU�K���j�FAF����+���}�!��k@¦�p��Ïz�!1w�!�ꎓ/o�����bԌ��H��̑�"1T�:���}���mз���s-F�����m.�Q��T�>��&�Z�2�s�����F��X�^�uD�c���sB���R�jH�7�&3.8�Wy.*		�=�3ĆG79÷��L2X��7R���[�� ܵBe�z�Q���d�ϥ�t�>L��fl�َ4����{���#��:�9�sffLc&���U��\�1r�sL��}�+��~��i�k}o�f����^�/�k��1=	o���F}{���D�?1F�O��>�2��d�d4>K��է�G�t ���օ
TyжA�޴sum:��c)e��K;&��;�To��_t%Q��϶h�^����+���/�e�_|��ƈJP��ӒSn}-�JjC(�L�C�г>%����2�C!0�4��+�#M�0�F��D�Ԏ۪�R"���epf,*~=����\�_��'�\h��
���|b۳]��7i��n����^��#џ��\�<����.:�K1P��		��$���E���ǔĽ�0��O���,�$�|���8�rp�BD[ϯ�)m2Y�n�n<gV����l�f�a<X˕c�����Jpx��˫�6��x�Y�1MU�s0[�W+����6���Ѭ��Uç'�8�Q��42Rp� �:dy��D=�ۉ�䰓�ʭ{b�����`�N��xʧ��4�񥂃���,q,�Bcp�� h����Š_��)���Et5�m9Fk���d�0�O�ZvA3D ��[p�f��,����t�s ���"��T �D�h���t
Ǌ�y�`�5�����w�_z?H�����O_�����m�����O����Ya^���(w9�Q�yi�(�̚���>ܡlG.GT9B��hm���G�}����T!��N5k!��) I5���zyc�m?E����ߏ�3�\"���ߵa�K[�#��	?�
)�i�g ;Zݦ�F�?�T�������~��t���0p	=8ܟ�5o��_�2-j'^�����'��P���,�"wFbTN���N\d�\���jz3 �:\GA�(��'ʸ	?����׵~Һy��������W�����W�Hᰒ��%�nQ��n���z&*�6�/���jF�5����~���L����A��`F�t0�0�g��7WI����>u��E�#Rh�r��?>� �JC��S�����L��J��t7�YA�یo��q�s���4d
=��޳Q���'������u����l�k�R�x��ӟ������(�h<��V�M]���6�xQXVM���[�d��'��|����z���m�/���ۢEN�'um�����9���W��8��ͭc�`b�>C����(����sY.����|(NFB��)�Ԡ��)�� �휏��qJ�� �O-Ϥ��{�eQ��j�S_��d�v��ќ�3�)u<�z����`���1Z��˱3_6���*O�+���������NM��3>�,2Ӛ8hĒ[-��S?���ȟ&�$`	����^�y�R�����.>|����n<��b�`�¢Z�i��DGz����LE��h�K<e,���Ie	|~X(^�Q�1�+cYr��4'�LO����~LxY<nP�����2� �wf켊5��{Z�1���z����s����B��Ӆ��{QO�}����}�	E�L�r�Bw�()��^��:���8����Y��!�X�A�g?�ÿ�u��_kxD�7�r�E���3�v��nQ�����Wo����_������Ē�- D�9��~���wW}N�	�)�ݦ0���n/A@��e�&�u;�RNp*W��V@��A/�m%a�����\���{�����q^�)�p��V�{��;|��p��#���҉A}�ϯu|��~p�1ye{�Y�O\O�?F�u#л�3FN�A�J7�7�5�Yv�֪ͨu�з*tNI}Z��
�h�������!���>mP��dZQ��U`
��6 1��u����>��6��k����S�������S�����D���8�d��a2M���?��?�]�=h��e�f�ҷO�nW4~�OO'�j�N�q���u�9ꆏw�O�V�2d�Rh��>k5��(ȝlM]������ez�!S�A~b;�Wύ5���C���ʇ�fOonP�<ɖz�v� ��^$7���.qT����a�"�/~g?Ɨ�h�h��rk���H�9����C��';�A���	`&֏auHv��!�g=��j�3nQ�PP8t8`|x�PLul���IA�!����kw�v��;���@1\�՛6�,Ū?kn�I���e%9�4�0��:��;�(���٢�������ޣ4������/���#�.��9�l{*?�+��=G��N����a�#	g0Ϸ�,u_�X�z�����寋"�zxt��<�8z���G�)8y*ѧU������S�Ǳ�)&G��p6{���Of�b���������|��ڤ/�7X'|<]1(G���� ��xD�9� 4\�O��6t�T8���7��r���7�8'8��M?-�x+L������،#�ǽL�����cO�7N;@���	��l��|���(s�38�� c�ic���M��fG���q�/�����;������>�y%ƶ�H�P��0	�� 
�ʞ���n��$�6�#�ȀA��f�c$�\TW�Us�e�r�`1e�%�\ny�����B/^|��=�lMW���T-.'8tQJn�56&�:p�3"�]�?6.ˍt��D<0���m��2`t(;�7r����K�g=�f��[Ү/�M�k�k��A��kQ�WJ>�.�p���=�����R��ߗ�rsʺE���:�&�`��xڳEn��>VzV���qs0��\7�c��0?�Vvz�#Qz��~��SV$̑����.�Z�ٮSά��� ��NQ��ی��Y�4xZ�us��7�
��-�Ҝt���R~!�)ϝ�1K�\�������^a����lhR�Lu�~�����^`�Y��+��<	Gr���C�����.r~��!QZ6K���d�k�m�9��ZI��-
zo���W �c�U4勹�4!T�sVk��O�A@�f ��@.��(��'��a<F[0��J���>&0ΘS����G��O���_xث}e��ג��R�[ki0��Fˍr�źb�ѻ<g�kp+���^F���ჾ�L=��Z���H�^l�ۋNDL�okYnA��1#X�	��l�����>Z���ZT���l��wX��[�c���~�3���G_?��P:R(j���4\y�p�b=�����w��:÷��Ř�� ��gc6^�G�Y����"�@����w��6��<]��\�y�i�Q��4��S岏�<r����Mj��#�j]�������E�w�*�#��uO��Fwu�QV�g�5v���5؜��6�ea��D�x|��>������FMJ��E�6t�~p ��?��k�������˿,���ſ���s/[����۩C��CАZ�*I�b�FGC|a.����6ùmܰ���g?'�4� �F]�>���1v�iRFJ��@���2���g�Qwf�1����#����>M����s>=�݋{Z@D!�7ew� �L8����vrw�^Uќ�������D|��c���Q������M&}�_��ʙ�5��Z��n�#��t��v�|r�H���-�My���Ku���ܽ���Q������Ǌ�~��
>��� �4>h@��0���M�.��2�\�ݏQs���8������'��PR��8F(�a�Rt�i��^VCG��h�˱q`@��JE'�<���	�E t.�}н1�1,ڂ-����/U_�]���Ϋ(
���O�}�a�SA�����7`������=���Ԫ�Ȭk�&:�o܁���;���y��rh�o��O��M9E��1J�Lh�uưʗ�\8�<U�NG�n>��;E��o�Ok�Gg����S�S��{ ��i:ï��I��W��WE��u�8k���'}dzp�����gS��y߭�\��Κ�h�q������y[l[-{�@����<^^�]���Hg��A�B�m���׍��m�aJY94��9Q��O���mb�����@92�fy�r�ZF-�^��*�2�����wxM-��"��g�P�i�	�5�V=߬G�<��(f�>k�2�w���<CM��EC�4ǘ����C+I9A�9�[��A�'�vk&�:�e�k�/�,bk���$�|@��ge�r�/{��[u�K?��E���x̹D�Hx��03���n.mO�8����l('0��hKg'hL��56��cX��f��K�����X��Ft�XsiPp�D�g�':FO-1�}�����"�)"�E=�1& ����"l�7�B�ǵV
	
�#�4h�yjӵ<�������i861�܉K�Z�jT�1U��Y!���B�I�Qse7���2'��PKF ���kx!�������0$t���_j��wRa�	7����[���Y���[s�̠d�����,(����ßTi
�\��z���R�p���XN������'��x�/G�*�HA�d�5EK�Q�O3x�{Ȉ����5.߂�]c2{-@؊��H��Oc&�2"�t�Bpx�%��b��ҳ�ps���
ZO @��BD1�A?})xk٪燖��{;��i���˃Ѻ��9-Jk��e+�����/b����q]$z?�,�u]�u5U7���d`A�~�+!�e�r�t9�/>�j�;c��E 	��K��1>>���iL�&Ǉꁁ��f'���p�Ha��o{�����Adf�%�vA� ���CoF_T�+Rz�|�#K�O?�E��8�����y�yj%Ĕl�	hЬ�� )|�ѯ1�a\Zʍ��%���Z��+R�3c��2���G�U�DE���?L��:X��&���d7(8kmBஏ׫�gB�G�x<3[r#����?�zש�����YƖ�ֿ�O�?^u�,��!���]w�D��O�-�ƻ��<���S�3PחC��m��{�{auϪ�����N��[�F�=���H  @ IDAT\M����ֽMiZ���}x�w9���a8ywo�g �P�w��l�k�}?��io����q
R��/=_"��;u�8�wP�^43�q�r:��1zz��g��ʔ�S��uW�q��6�nw[�i��,f�if3�w��ų��V�o��u]�ӳ�?r��'g<��0|2��M���,���\v���n�O��V
��Kp:������߽�9\Ѥa���������-���k#9Ф�h�5녣�1��\��*塄Y�m�{��+]_6�RDM ��6��4�wՉp-�4b���.}��8J��r}�S��o���ʀtc�W�� 
�j���۲}|�ou��W-��I�p�^�k���}hʾP9����L�O�Q��v
��1?�d%�_=S䀜��C U�)�9�.���*���TQ��o��-��3H:�r��+ړ�n�����y_6J�S�蒹�>�Y��M���EQGĜTȊ�v�i����Qq��ހF6��|^djA���P���Wf���a�o;/��昆�ӻC���e,d��Z=�B����Vw���z��5�^�0�C⢋3�9ě�^K������rZ�1�<\��"����Zׁ�t��(���o2��z�4��V���!X��M��A������yvуi �m̓����O_����VEyQ���7�|��?��Y	�=$G8�v|[�D[�z7��Hx,(}�B�?fW�}��ʃ7��&�wsP��������w��.���z��)@��١�J�D�ݻ\'D����	��3]uʐ@'<^��Y)!�_�/���Ṡ�!�Iؕ�0k9S�s�@���0��c�&��ӥ���{4�}��O�x�9Qyn:lW֟�$�]=���? �N����ғ�Zg������Q_���Zi�	���tL���ꗕ���T�5j�k�HL2eَ���U_Wɸ���u;jC?�uI�1�A�๊���J4�]Y�������g�� :SU�[��TV��Z>�sz�>Yv1�oF>�S�u�qr������?Ɋ<�x���P><��n�����D�D�t�x�n,�n	��^������W�_��_����˿}�o~�ŋ_����),�}�G�L?�#���F�U_��W=�)�		�g_��\��>؋���Leݑ/OY��B���p�}�e��?��2���l�>?�GJ��UA��������6���z!�m�^�д �Z,��]�/��)��^g]�0=�~g(	�Rs��ftwo�R)���_c2�@��ɬǅ��(�"�p�[{[�#���W�[�qTʫ���n�g� �o��Q�����|8��o,#7�ҽ�]�H�(�����6e'��r'WF�����y��[�2�n�� ��dw`��ykV(������O�D ����+o��:�7^J��hEK�jR�G�<!Q\{"t�8)�r:����tm ��§E��;�tQ�Vο��p�&��g�/љ���s���`O�y��w��N7kVW�uё?GD��!YQ�t���L�/�/��q[�2�ϔ���c�KÚk�������zmC��P$J�H��L]��5�`yz�գy�<"�)�r-��<w��2���pe���x�(�g@}!���!�d����IH���q��w�W7���F�	#�pt�:���Z��TP9��Z+��.fZ�Ia-�__�<�N�m3
�:O~��s�,7�Dl4K30��y��c5����>��Q,�_N�*�2S���+V�;���ڽ[u����5���xs�%��{$�����S�{���P�:��W	�3��d�����5�A.�^��`[�۾�9�9����A*}��5As0C��^WF�~�[�$:*�s�K�343�4N/3[�7��O��&��d�0?:��Y�g����W�|��?zCxIG�`>�?�/��^y��ȝ�_�=�����	��=��{���9���0H�����^/^���+�/����7�fo�I��<��Thcܼyn�dʅY���ۺ�	V�#�>�z/�����[���<�8��v{f���!А��cze�sD���ݵ�o̎����K6' ����(�8�A�8��=�?U�g�5E�������p�������}Hyb�M�&ɂ�g�.<�����8��s���i�ѫ;đ��3��'࣡L��7M�ђ!�ȫ���kn^B�rB�)��qVϓ������jiQB�?�(E Z9�cХ\F奪����6��6F̙>�8��������-@c���pi�P��S�ꖿ�s����7'���E��`�������떤�۬� {`Qԫ׿>WR��{�`���L�]8��Y7ǿ���2|7�q-64�p-�g_���s�0ђGC�ES��W�а�A뿵H.v�ܘ6�|I:`�`���Wt�ބ'r��G/U^�'�)�/���V2?�!bc(�(yp��P̐��)(#7fP���B�Z��ǧ,���Ǵ�)�R����gˤbJ�M��s:��甄��)�_=�¬5�\YAa]¹�Q=>����{��"�h�n5G��E41_2�t"M�f�<|�֝Li���\�X?s��L�/��=��I��J]S�5)����>j<��P���w+�n���mġ�R�S����i��W�������}��n�^4���C��dV���� g�5
p#7����f�Q���݄��&|�0���আ
:�60nZ����|����i�E!�>�r��~��=���G��S����|�DTv������K�.X8���ӧ7C�a�vKߣ�cs�oPTtRuۗC��[������O�&�)�gOq�a�Ixs�ץ���Ho��\J�y���x:�������JgBL�*����=O)�m������/�ſ�W/���2��fL3҄�pN�N	���t�-ͣ��ҝ'�-���F)�VV�\�@u{ʍ�ʣ��/C술.!��{-g�7�\Jـ�-�P���B�w��~�;+�xܛ�j��n�/6�ጕ�����pf�i�)�29��Z��2�^�1�L�W�	>>ީ���·�fy��Ǵ�!㭌��k]���L�c���jMɰ�XP?�ɘ��4��	�GWp�оp�X�w4t����[Q5��{Թ�)y�t��u�9�9 �P<8�C��d��}�M�ú���EA�8������IMf��DǺ{n:������\uЏ<���$�	+���3ح%�c�͛����y�F������w����,��a4��V����_-��V»�jO�v�?����3�����I�N�M4�}?u��IӐ�t��l���W���U���������U>��8�d�xa���[ҧ[��d��l���݈�?O<|�Ǻq�PVH%�[	=�N���нu��|�B_KC��?n���t�?�BA�#Fx
6E�A_��Vf̩� X�`�/E���a}�*F�wf`H�k�Q
4) �|�x�1<X� ��p-��rx�2y���2�aSbP��� �0r������pGs�<PS?������k�Z��G�x��)q-G�L���T==�1�i�@�����E�-��,�(5m���B�sPx�bx� ����Vt$�?��u�	G���#+�@.�Z}ʤ�q�L{��YNE�_};t>s-�,j����Э���΀��F6���s��A�ϯp���36�Kd<�	)�t�K�$�N?Y.|�L������߽�}Y~�Q�{X������p���t�7H]�����s����!7��ӥ��uS�w�Z��mD_4ȄA4��<4֧�a�;���Ҽf荁G8�φ�2b��PV�=1�e-��7���?)׌���wʅ)��sƢ��l0i]�`���Ypλ/�H"�x�4&�}��v]����	7�z�B<a<B������FZ�)����Zą��N%E5V�k;S
|<C���y�;�D5�n����9��� ����ĉρ�3��r�ѽ.���ᢴʏ��\��qX�	|^�?�j�r�͒C8l�B��c�iJ���׊>*��@Ti����T�Zy��-�Gr{�p1�}���9K��+2�W���Ѕ���!��q!ᕯo|��ہ��x����W�36�z�Lt���SE�c�:�278[�*��pQ�+�Z����7ץ*���W{�HV�;$��������������턹*\7#=�X�ʝm��ϩ�OX������N9��ZǠV	�{���ЦH��Yy�cl�d�IR�0�zK[�Y���p�v�7$ *QriwQ�\)ܞ�A�]p��2�=�4v�m��5��`˾�e�����,���G��\0x����1'�B/g�!-�ǳ��
�iMB�����������؇؏I�˱���9<u��Z9Js�+>=�Ol_ 2����g��G�7%�}+��<N�ZA�?t'?N���Q�������!���}ך]�co�DM@F�#@�3Ρ��c-f�Ϲ�']��ˣ����pMW�a����Xef�����sN��3���΅Ǧ�B��z&{| V��w�ߕ�IZ ��t��c����5B�szE����֍�Z���ސw�<!~?�����`����듍��8�s�������׈8]P�..����΂��0m�Dk�����y�{թ3F�#��$��"ĸ���λR��>胲��̣����1n� j��>8�Π<���$ ��DᷟÏ����
_}QJ�ow��[����}����9t�1f���R�{ǉ������$��؈�,z�
�C����������р1x����_���]ӱh�0�����f��"<rEN�>\Lh+��U� K��ko�4�F[�g���*^��h���D�P��2\ˎ�������Wb�0��0^vx��O������2������6ޕ_ZD�KӃp�<Y/�E��p�{��X��7�!1�_��L}��Ӟѳ�+7��W�bG/����!b*��0����] �./��� �|�D][�)B,��)��,h��e�����~�ۜK��c���xǒAV ���9Ҍ]��;YxP"��w��^8�� qo�:6</�qj���~�U?(x��*�H֪���\��:��	)E-�CV�@���ʇ�����(x����_�}5?C:��N	��px׍���'�p�+��ޙ}~'��F�#��㪏^����P�nV%�-�.��I���acN�=H�^�>�p���A�b�}ƶL�7��I��a�VVO���,j%֚���q��G]�$?�r��!4��$g����o��ܖ(k����sp8J-��V*�@��Zz�3O��?m�sb��m3�"0'�='�Խϵ��r��ú=��t���c��?ڝF�n�`�G���~W6��i4�t�w�� �����;/�uB�T7�����R��a����j�u����DX�]~�'Ly��g��q�ޤ����Ԙ�յ�	��D@i���[>�݀~�]��bQK������������?��?_a(��U�V�ƴ����������E�-�)y�o�	��{;�W�Sum�9!�6�D)1
sOI�W B��?����;�ʉQ&�����b�� 3>��<e�7��)�V3v��x����"X�W����&{���W�>�1��ON����s�e�1&X�LA+�n>!� B~���|�� ����)h-�����f>��0���rrk�Y�JN��`��C7%)���Q��ByNv�G?�Nx���-a>DOT!�{-��co3^��:�=Gx<��U���Z֪ ���3mg�?;����E �_��G�;�!J�[D����#ju.���{�^��rd�	'G�;	�/8>��El��V��7�g{��z&G�C<�N�_�9�A�?�o�Tm���V<}����2|М��@v��W�O����YB��N���Q� �v������RX[��:x��9f���祀����l�|ֶ3�jb̯�Ǵ�[U�Y��޾|]������W�$Sij��qs١jz��)��o��G��p3	#�)'�5Ԫ0���4u?�]�㘕����N��]}��V��9�~�ĭ���<ӣN�0׵���/BF�#�Є��m�س|�O#��[t�B+�?���M.�{j�ʟ!i�����ue�a#���}���27�4]����g|���u���.%���ݜ問,�_��P���G�4ϳ�e���Ɂ��*�ۨ{�o�%�k;�թ������ᥱG�o����֟�N�dy~_l���u�,=Mr R"@��w�z���f�]U�ǒ�~~�=2f���~�ٱ�۱�Zz�Dќ�6'Wᓎ�J����!5>�܊
N�p�Nz���%'�n#����(�W]�"�_��Ά�{T��
�l��|8	z}:� ?��>�b�5��wB|z�o����#ܯ��e�iT|�
j��%X@�|l�ٌ�6�m3
�X�Jb;�험�(��4O�7��`�N ��ȃo��w'`���?ofv�[�4Z%O�C1|��P��� ��-̝��g�(�γl<]n�]�=��~��O%�K����=�<G� �[���������~���+����1����l#������U܍UĢ����O.
���.|R9�'��S�诿J	���s0�dPh>5�Og���z ?`�oS���]���Uoua�7�ޱs��ޕ����#x^������hx�T�����;��Ɩ�9�wu3�9�k��f��3�#�cl6����e�-�:Hz3S�=��T�U���G$P���'/�q�U�!�%�F�t���`���~�틿��/P�XX���n'�T�[�彣�e�D�-�Nv��$4=S� ��4�û�p�̣l�{ʷ���ş��/�� a���5J;]Q�t��Ȑ��o�P�oyS�?#���t��0b�Z�e��^mU��g~�I?5>ȨZ�$���j���o���_�w���Ɔ��xFk���R٧p�b��r	f��+�����w�?{#���9�ƀǠĨ
1��&�d�`?�����:����.��vhdp�Wҏ��Y7f=Ң�~O��W�s(��2�ƀ�8'7R��M"����|�<�_�㑾8<�����,^s�A�����V�Q�Yw�h9Y��`�L�zr&�B���+�H���h�?�`㌻�%S���w�m�xI��n�ӽ>�������I��'�iYi�9�Pl��Ś������W4"7 ��K�e��{�Z8a����v��Џ��̦:��D�!��l\&����@o��T���������j��ot}w"~�Za&������i�f�Ǽ]�9�3k��S��f$��/�@��Q��%<�����l��3A@`J��t�����z��+f�L��3 �����7`�`}�.����z�Ze�G��5+�e�	+]���{ҽ���X<<�89٫�s�)�R>����7D?�F{�- ��Z�LB�)'�*��@��wM�.8�rt��R}V�>�+O�[�w��g�`�ѿ�F0�	.�b�F�b��q���(=����bP��c�S��
V�ɴg���z���+��̩jӷxdW��V7��q�����[8ݜC�B���ᚁ�?�`Z�m�#	Μ*<f���a	���?i��.��Iҭ�Z���[Z�k�ԙ�����C z9�?�?���W���l^�����yc��F��#�hc�Y���WJ�����K[IY_��a�����Ӌ?�c/�)����ƅ��&�\�k�t�L��Y��M��_*BmHR�=�p���qd�@^N��iQ������,E@$�����@�X߰>*/��H�n���>STnc+C�x�c\F"��Z��cG�Q����i�� ,
q-�
�y�\X_��	��0�ȋ��	M�1��+cJ�JoL��2TŌ-	�7��,��M�Ö${k�z�-8.[�+�P��������r
���1]hS�W��<���n��р�K����f�:Lw��d�����d�GfZ�����V/���^|�{�k�b�tu��Ts�9.	�p �זco�9î��[r�Һ4��d&�:>������M����*EO��~M�g`=7��v���	J?½F�*�ӭ�vz-�P�qlh8�~�{�����4������r�P��O�$r�V�OuO~���u��jD����*<��y�?��O9�C�KD�P5d�*I	ϔP�U&/���IW�)A���ی��r|jJh�N�����T�yZФ1pקlO���^�S�X[�C�F��`�a��bk���U#����'hp/�\k^b����)����_ye��mB�׾�w�N���>ge��;��QdNhא�� \���?"��Y�N��s�Lʢ��z���7}��4e0N��?�/�sjv
��&�94�6���5%8�I���T]W`r��W2#b=0���p�����}M����*F9�Q��������y��];�}�6�� ��V���/����o�-l�$ޠ$z�:�_����̔���3���K�G'��۸�Ç7���+-`,i���Ur�{��=rݲ�����}#��6/�1�f6��}z8�g�3T�o�T���jp�QV7�>o�+�nҀ-�[�_t	���y����:y�}�5�Ta��\���'^N��"]��X�MX6�$�~Wc��E�1�j��)V��LG�!t\-�<j�����iE�̻Sj/��U��;Eh���wJ��݋��A����Ҝ�ڢ�3������mH�tNgϺ�ᣗrD����t��QQ�����3yo�&T�3e�Í���+��]>�R�=��A�����:�Ze�k�mױ�@&x�7z�O��O�!��EaE"������
�9�w�Z>d����oN7�8��u�p1���� {�ƺw��w�<؜ȫ�l�Ch��NE�]=��@4{{�8���_��-Y���	�N����D��iȻ����g��H������,E�8]J�p�4���!��E���9ݶ)j�_�OtҳM�vOT�+��O	�i�T=����|��.��������+��o����	Ǩ�~mz���a�9���gӴx�}U�`��ry��3��B�>��V�k�7�1f2���(iK<Y�ʭ �r_0ʵ%�.�G^e)��6¶����R��`��@9�b���2sd\mC���dZ�g�\$�(�������ΐF�9F/��.��<���2�}^�3G���I�#�����y�3�U�V��]:C�'�ӿߞ��a�gX�)j�i�����s����j�Y�2\𫫻'�(�?��`7����.�o)�p�g8������W]�ZA!����f0&��6�hPy��5�������f�C~�tN�N�� ��"�u�:C�ˁ6#WAzJ���4����ޅ�����⊂^�����p\��-��� 1d�����1�P�<�Y�3�s"�eg?7�A��x��$�Js�F>0n�t;\�v��`=݃E���~���>z>�Q�n�![��,�yȾ��q�\	��R}��_������V�HA��S�!�S�`S��Ԙ$^��n����R�q?��;	��k� ������)���Q./���.|"��nky�"%�G��9��d�0]�Ro �7���Z�7���nh��"�#��r,��EcƨLB�#SY�Q�O	a�%����dRZ��+�M���®�����_�E9s��9�i L�������['OH5�^���X�<{6�K;��0 p��~���Z�ӏ�����7,�7-s v��f�ɍ^�7>jt�F�~�A8��3L3�Hᴴ�zқ�*oV�f���|$� �j�B���=�<6��sN3���`�V � >�'�Gr�1�D�t�>�X�:�&[f�e���⍣�[Q�0M��(ϴƐ��ޢ-y�O�c��䳌Ԧ���*��[�QH�U�M�#�~�s�6E������A��T�������ߎ����9�y�o�.&|]�6si���N����JbC���Q���#!� ���;a0�-/%[�	������:(��HU۪������]}Ȓ<��`m ��pR�1�B��3��/�)l=�s��f�>��LXt]�`�GP'Ʀ��N)��6�OC�w|6z���pA0�����.%8�[��%|���_Ւ��@qV?�{��:Z��o΀Y��)���Z��~��8�.ۃ�U#�#8��	���1/bZ��^��1��{�0��1�dt�q9G�����ßcIk��*|�����A�R2�e3���C�	������a��#�mZ��s">A�/j��y2�fN7����fZD��i��{���$i\ߴ��̖����Ʀ6~Ň�c��m���7��ƨ -��_���5]�F�8�Nj�ӛGCK�8֬��TS�w N��#R���V6��~�j�P��֨�5A�c��A^�����v��!t��3����G���C��%�{n��k��6D�`���KZ"Bx������O�EȻ2Y�B�MǤƅS�E�Z�,����)PH<[��v^��J�S�S�2`���҇�6���2Au�5\7 ������	}:�:��1��c~��2�W��*�#���"���j��;�=x-Z�$��Oi]�V�޽�j�{�Z����8'v��jE>|�!��Q8��GD���ͮ����L����Ԕ_�GVN���#�A��1_4(%����M���nts
�r<���$���2/9�ʍ��=�L箱�6 �TP��`v�x��x���x=ُ�3�E8ɁD�D~'��b ��Y:Z�N[l^"�a-�Z|g,��P������0��˞ql��_ܝSR��_��1�"c����Ҡ�)v�$�ET��/餺�1����K��_ۥ��q��Q����L2R����&��%NC4�9�~�Cvbc�>!�	��Ɩ�R��v�iPZ�'�cRf�9���S�[�˸S:�~�a7(&�Yز��`�g�?��i���3���+�$c����'�7=�����P�t����T#��$����+��D�K�?��L�����x4���\�����gv�}ݑ�����[�~(O�~�Ύ�Z�Ɩ��3�����8
T��S�e\�D�f!���$���<�2zs�S�d3.C�g;j?޾����׌[���C/v8ˣ���&�M����#�5]I����E�����^d����dB��s&��o��e���?�Q��K+���~w�0�gr�H��[_"z�����|g?Lú[��"��?GL����"�V�n\$�d�[A��v4yiJ�^�I0�;��L�8Sg|i��Z�P���Տ7�{#���
�6E�F{!�
S�c�o�[�"���%��<Z�L�4�N�4nf����י�o$6"qQ+5�Z��S�{w�:dŏgZ�у<��GJ���;\��m��{�/���|�����7��CY�w��_:[��=_��#���Ev���8���%�nUy8��^��ĸ�aLJ�pZz<g|�t�GkY��]���n)�����x�2��x8 �c����u'�^W�\�Rި�~WnJY~<������7u[HrJYs,���:r}�����u�tg��3k?To�" HD��e+��(G�X��٭%�w|�q����+|��+ȓ$C�LQ�[ӯ�%��ee�Uo �~p���(�ǎ������,R����O��4��e�+�Ɇ�.g�����np����I�#�T�J�j�C���دq���h��������Vܱo����>ġ���J��t�s��͉��կ�(ޗ}�����y��i�[�<DD\�=��{<{�cN�� ��o<�Ɯ�(�wBX�CȌBZ��F�OAk1J7VR����<���_��B�p�'�b�0X�e���
{��_9�ߞ�aB�z����3����_k�q|V^uU��9�>��k�*� �>�cף���)�3yÚT��ae��7\�!l�L0�8���]�k�rPxբ��G��w�;���U����T���i�0e(��i}��$b��j3����x<-��8�O]�#���>'�q�8���N��,݌O��t� �k��Q`hO.L;�܌Xy�ZklK�����t�y��9=e���zս%�����,�l`��ݘM���?�_�r���t2zY+Қ3��Mt��zƖ��_4H h���@b�6���Lңc��B���J�o:��C4�V?l�Z��"Qj�[�V{z�D��������s�/�Fī��ӽܓ�L�s������n���p#wJt�� �*2.�:z@���2jʘp����XdQevu�m��S�C޵�Q쫑�5� ���|�V_ �ׯ'<�@�fȻ�?�W�Q�����q,�E�_�G`��~
g �n�Om���o�TH�����p��R*;x�m�P2�/_+�俨n\�2�M%v��6%�R�� p$���>��d����WY����}-��gn�j��M�F�צ������"��Zw�C�5e~��e��V?�DrZ��*��`]R\��讁�$28�/�%e㷴5/����T��fO9I�����ݲ�Z���rtᨾlĠ������a ��ij��]��G'���D�R�;���q����_�+�?�n� x۽1u�c�Y �Iy0VȺi��a&?��
"���4Š�5	�P�V%��b!�Z�~#*5��M��w�x��ff���[��~�b�	���	:�g���=^3���w�}h�6�9,8��a�y�����WY�,��>�h7 n����Fu��=Mzݧ���_)�dU"l$�'��{=����G? ����Պ�Rއc���o�a)����rʥϧ���Ǘ������3�T�4������5�1E��ѭ >�%�.#<w�9g��>� g�CO���&�V�[t�҃90;}9a��
�Y��T�9�䍏����)ץ����h�����t��2�g���zf�p�����������Kp����E��/�p�Q����-=��{]�5HHi1�Jwh�:+�5{]�ݟ�":6ek�Fɀ/+��s$��{��2�߷�L��&fOy�(��UeS�.J��Q��<>s�>d��7��+�s3(���J2�I��Z�T�Я�dZ��Ӯ�ߋH,^�Q��������$/�SΘ� �,��G�;r�򛦚x>9X���L����h0�~���`#��>|k�C0��+�A��������V�?�T��5�Ɂ��͉x�c����<�]$VK��30߀�o0�
��:M�}�˝�/�0��9��y�	����6�q�S��n�u���7��i-j4I�Y}[���I���^�N�\�co�ΑД�.���0;@Kׂ�p��Ǐ��Q%��[=%�+�G�=�~ûRˋ��n�w�rƛ�I]�R�GN���y�L.���Ej�5h�٫��K�6��mʔ�����S�*�lм}<����w���R�ٚ�vP�sU���HK���j�u�itZPs�p�J�*�J2,L�w�7���y��������Άc �S��:.�UE�s�
��Ƣ���Op��p�s|8�Rg07�g�3���m�ko!��Q]����ni�D�~$��� Ӭ��@�m����Z�E�6�����]z8�y��#/~�Fݫ�B�
W�	_?6���L�N��՟wЮ�o;	�He��`�Oy�}	xN����I�qG�˷u�'x`��*4Ytdc���7gBau�Rd-_�~��g��[wA�)���τV�V��>��!k�*8҉.t%�ւ&}p� :�!���]o�j�"��z��1=e
O��d�_���)4v��,�;�{�:�s��y�&��n�����V�/��ZW��v��C�������$��"��)|n9��=1��9 >�a�o�yXD�y�yݷ`�w�����C�g3J�n'�S�$V���Cݸc|6�˹����?�q�W����^����E��P1߉�k3NB��|�d����������v<��nL( �x\" �`�����X�l������u�/��y�PR���0���֎��%Ha����I��'�g�{�y?�����p
��ԿG����½�i�i-�`�thx.z��\KzZ�F����ѫ�9�gp���<J���op�~�T��{6�t	׻��R��-���`�����A��c��dĸ*A�clҪ�֗q�gP��Z�M����� ��O����A���Jp�㕌�rϻ�n��s���2���1�{�C���(���ױ���iY5#�u�bM����9*�*9R��O-T��.8X��®���[:4�~�2|zUor0����n�?��on�_��O����2�7?׭�g�	?�U���a�4產�N���=�&��s-���������_�H�Å)�!ͣ@\¤�[��z<��N`����"���W���)P�����83����I �Om�(Bd7,��[��e���	������n�O �w?z|�U���Ӌ�F�9	��Z�e��c�0<�<�����>������9��}
o��3��dj��B�)B���U�F�ï<�������{8�;u��=ɑ]^Ƶ̻?^��9"��*�(��m����#
?��e�Br"��3�o�������,�e��ח�N|��ŀ�RtpH�N2��h��ݺa�XPN��>�N�����ҁ.��ρXl��<�6;'Vh�����������W��z=�O6�v�v8�+~H���|#�/���-䄊j�������N/^>N�S��P�xN�%���G��a��c�D �ʈy���_��������{?��ub����쐨����A���S{��m���p�-����<GP�-]���W�dP��4V�.r8eZ�yKyҸ��r~1d4Da�B�������(�PQ����Z����<&�|YfNg��������v��n�?�u7�m#R�M�9ţ�>@%�<�rFe�9\S��e����սɰ�uo���{S�ɠ�_�@)݂9�?��׌�_Q��%��gp��4�w0�F�K.YNY�V/�v�{�]l �Yi��AD��&/pQ �3/r�.�(L���d2�偣O�����hٰ^[�Q������ $^��%���q����{��tDD?��W�Y��ԝJ�r��iP8o�4G�(� �9<���j��;M�u��3���x�o�b�?8*�v�V�є��T&���R�&�FOt��̋�M�~��� �P�.��__�����S(g��{d��0��^�1h����iyq�Y�9e�R�$l�F��h��-�Z�����'
˫�YS@�_W��kU��շ�[<�m�9�K�i�̮B��t+�_�+�3�]�X����N��wf�k�Ϻ(!�->��W��_
�~y
��H�Cj��#k�v������]_���;�i୨bK��
w�s��Gk|�g��Y���)z7H��g��w��Z���K�u2�9�ɚa�(/����fi�S��9Wa��M��P�4���/�k@�0��:^�Y�x����I�ۖ:��Y���0�۟�,8�m���6��8�ǲ���q�t�L�}y��٨���Eu)��|�!\� ��Z�~Lgv�6��Dvur��^��q&Q��	����q���?8�52!��'!�RV{��7{q0/� ���d�>N�$6���m4Cg�����X����:n�Og� @�*C�K�'��g#F`��@h!x��ܭ��oiL	;����<�6Rʓ_>y�$'��Sa'�U�8�&��ƥp��AA߼�pP)z�E���<Fm�kZ���Ts���X����	�)c�YR�o�e���ї���wk�"��rB\�Á�h�tuvEx5t�]���#��c�Э~򓿧�75c�֐|j)+H׀�MJ|��)T�l�It8��u�M)���Ӌ�RY'c���5��Q����hZk;�Q��� $�,?��]4��D5@���E��sO*˰�32���b�˝A����U2����L;���<�B�i�i��~:
_2;^�)ڐ'M*�%��Y�г���+bǅ�-�QV�C�o���;c���염�r���"�?D��J$�� �Y�_N+�_;=^=�q  @ IDATE�I���$x[#h7l�7��:�t{,*	wS.^��\��O������i����NH��D�a�+�P����3@$�G����������cR���}D Na2�� ��Tt��?�ߦh5�/>��z{XG�L!��`ޒ�N@N�m��sݫ�5�e�Sv�f�I�,��1�[����	7�9/c�+�@��>o`-���؀%�
���ǭ����Xy�3�~��f����s@�'�#*{ܭkS�s���-������q�ݦ\�0�ā���EG�7T���i��#�E�Z_��>PǇEC(� {��}.Z�+-5�fp�!�46|/G:�ި}�x@^�!�]���tT+��N�˸�#>�Ϗ��+�~)�c�m4������|���oz������O�Zr8�9���%���X�r�l�ry=<�}�{]��1��0ĨջU��MΉu�0�gTj��͏?����7�ԋs�����/Ǡ1+��%{TN�@	<��^���֌g�b�xs���R7�57��o�=���q$���{���Ϩ{�u�k~~��#�A�\�J���	��<�����)@?V�EK�:a݋�`x�	𖂑��v�g����Ts5�#jJ��\�i��S).����IK빐K�%��2��B�i$y`�#��U��U5Yj�&2Y<Zo"B����Q��1����?lM�A7�{������	�A���cXƜ8�u���}����'KN±�:������X�b���tq޽��A��>vUb�	��2<�]	Ǣ�Tp	.ۆ���lQCA��d�le��q��[Hv�@��]k� �g�k�����r�aoqW�䇧$�v�g���ܦ@����(�dl-�>�mP�1��.18F�Ï�R��w�l���"8߯�+�9�@������pΠ������~�Ak9iJi}��������� (B��2�cZ�ƀ��7��!�ٰ��b�<��ٝV
�A�a�'����C;�b,E�/[�7l��{�z��!ny�*����a]�_&�.ʨ/�ih�8s��k<�_�}�~*2x�G�"��O쾁��8�0����)w?N�P7��>,� X?"�̏B��r���+-,G~G�ǟ�v:R�� ҌP�|���$"09�P�H���aC�9��tB�{?��%���EI?�S�]r.Z���)��6�+4�ʟ����e����(;��`ey;)����}�)�t����~�����EϜO��zU\�3'���}P���׻ΰ\��ov�(�'�_��À����NN&�#�'"���{e����^����P�/����s�tf۹g���ձH��!�ux����]>i�?p�~k�ҷ :n��h�Q�!�0� wz�?��?�� F�^��ZF��U)ai��㑴ꁝ0yv�Z��.oA�
�F������W��"ΐF���>fȶ����_���)��,�����Fn����O�����Z��::xc$K�HNgx(�#��� f3`y����ޢ�-��>O���e��,�<�Đ��>[AXy���OZ��uq��R|tkY�$xwݤj�zc|����m{�r)�V�<k�кRr�JZ.x���������.ײ.��d�{|?�}�.g��|\�����ڬ_EO��w&�k<�=eF�$��m@:�����ΎON��n��P�aEk��ާd���F��`����7U��8�h����5�}X]���[��S�A��i@ƍ���lf��lIYn�Ҷ)<x��x��O7v¹L_�_��A�P��~��!}���y=��Sbds0��0�i5�^���`�Mg��[e�fIk����oo�� ��	nB,�)�,�������5É����)(z���C@�M �7�v����4F�D`��;Ah���"+	3P��8�W}_�c�t6K�/�
����1F�g{9������\��Cև2TO�5Ƿx�i���~�8�	��tR��DFb�#���x���x�nӝ�pNm�RZލ+kֺ2��VŽ���x���@ƕ�;T�9�c��4��s �<��MWA>�OQ���N��L�<
��:����+�Aa�Q�����7uM��
��j��s���U���|��Y��3��/ˋ��T\��~�\}�l��1ȓ�᧑�8����XS9Gb���e`�.:�A��{L�R�/qb/>�_�L��?�ǫ�����o�6֠+��ef����͕Խi���[���S���{򊷜�����_��[���V-<x2��}��껧���&q�W
Q)��$�nq��U�0�"���� ��}�[O����	��zSHDQ��0�;(�6kO(�9�30�y�sj���1lB���<%�d��4B�Έ��h9|�z�	6xm����LJJW߳EY�_R{MVeV�^��<���T�7�k�X���_��{bi���'�(�$�(�쳚�utC"�)`�~�`�������=�ϲ\4quCcc!}�����|��=�2ݹ>��{�t������Ȫ,K蒴�^,��C6�W�1�L>�������u�$z�H�k�?��\� �O>j4p�=1k��Vȗ�Qͳk�#���F	�Oy�'�h�k�y��a�R���5Ѫ���wXn�D���B�����h�(���y:م�y�z���F�#�B��������;�?@�3%��1�A�
��j����W�G�Mq���[�G�3i-��G\Ѝ7�{r=�zΠ��)��D��H\��@l_�Q�-:���<��Q�K�^K6%����&�O��/mD�{ޛ �y�Ƈ�7S�;-�B3���z�l��Bn��.�^_Q�Ժc�7߼[(?��0��;^��sBs�����p"��������+"���]�4dB�3Q/�?YM��_?���r�S��V�Uv3_⏿\{Fp���ڽ/�̱��=F"��_f��y̡F+�
���|4�Z��u�C�Ko[�����ߪAN�z��~�xp*�w��9����k������ä
�7����ƃ���������;S$��1���JH��������3e��!�L�s���}ӽ��xOV�������1�Z��Y�,z��|�L�(5`E��oz��?��Ż����i�<�)��oѧS&!�o)}^М�4&�I��JF �c|�X��k�Z�{#���x0�:�ь�3�͖q��8�o�01�)_��1�����;��b���'�N�OA�;�E	���л���K8���<������@U������3x7���:R�ӿ�D��Y�LOky~'��>�N	��TN.v�7��0�u��0���H�2�G�ޙ�)Bd�h~�%�+]�}���i���� ���㷢�^����{_�V��&�ZF]-����oZ���?�/�)�H�\M~�PZQ9�����"1���t"\�g|~���Ə�c�n���N��[�?�Ȣ�V���fn�H��������vSzkt��x���e�MTC�,Q��Qj��;��{���S.��7��Kt�[��|n�6���9�f����y����y��7����ӛj53z�>�$�S�)��\���O�͑�>�xE��)��=��_�W��砟<k��Q&D��f��qE)A��n�f�'1�%4U�NS?��!J�={��]L���Ar�ؠ�]�Ko�+f�mBg�Y+]z��,���9���O�5�(�a=}�7#����W�rHBL�R��e����IL�wG��������Xǯ<�i���'_�yS��|(�e	�)�S)H�Z��'����-�ܘ� ]�4�`a�Z����Kh��5xq��N����8��q�Y��[$��2�x;�����xex�-��V��VQ�U�f\��[~O��Νq4ճ�T)���VpP1qF�68����UVt�n�E<7�	�r���3Y>n�e#I�� ���2��8��R��%�M��|��o:�����o�}�׿�.>��� �g#�VWm}9���\6��E:U&�v�����u5�! �Ѹ,��#�%kL���[S�����ʁx%��o~��e�=0���n��P�g��P.1�>��^��b�2�-։���AR0SgS��mV褐�xc!)�����Ro� S�~>0a|h3��@���>Z=[��3у����H�Cͮ'��z�l�(�q&��v��A�������/��'�"�VU^ol��⣽���Wo0U��\�76@>B�[Sr�"ͪ�R>�[+��3g�B�(W.����7:�#у��oq������cE%�~;���lk�\.f��a�2�=:\��?u��tuG�s�������ׂ�Stl�F:���9�7�'m�7zD<յ7m%������a� ��i�H}�CnA_tQq�ߧ
'Sy��_���;�5rx�CyS�f�uL��}� ���}��?���F�	p�:H�x
�V���)�hU��0�)���d�������b�ZK��ϑ��H�3Z���W~a�h����Gxm�E8�[+�1}��U�b޼'ϲ�7L9�ȆC�ܕ�#���N�d�L+A1���lt��1f�Z��/P�Z�o����HMs���q���=�	�2X��`��8�&vOiʃ�3�GkPg���3�U%�=x��:���i9��Si:c)5z�R+���8�zӦѦ�2o�B�l�6{dt��l��9��n����9U
�آ��^+�6�F[�b}�Թ2�Z��l���w�o~��dvAi�dk���cBs:=�@���\4�x�E�+|�}�m��S����;'�9D�x�PA�� �a#��N��c`F�oG����a�ـ�aS�w7��֣�[��U�+r��`	�t��%8����-_��Ai���~�A�X�~uK���@fG��n�һw�� )�DRMX�s�ll�[�),AY�H��ן���=��������*�z��zqwlJxJ|u:�\�0E�et�(0%5VB���Y��e�������Sh�^5�p�ϸ83ぱ�eX�Ńy^�9�a��*�Z�Jb�<��U>g���=<�Q�S�`��s���?�Eu����l*K�������l@��6��A}År���d��ۺ
��|�<�E,sr�7����p,/��nWa�uʉ�e"gy]��)�C�(1���ڀ�+E`�"�` ���AF�A��ڱ,ux[+����}XW�\�_]���x;rOz�q���-dEp�0DW�s�h�7g�}�-�f�~-�u���A��clǐ�H���@��'��p�K�ЪxF]�&Q�o8��6��W|����z(ۍ_Ź~�](��U��EU߼�]�|�L)�͔������~|�����ص��PݧH��B"�0(B�
��Ӟ�猣[S�?���җ}&7�#}v��3�nz���s��@��6s^���|s��$��)_΁�� є�'�3 Lb,�p7+�⇁��>Ä��BV�%�P�Z�7���'܍�F;$�mq����?Fe��=ؔ�? \\����:� ^R(�d�xD�����]��}<���|�-�h��a�R�c�?�\���P'�@���
W�x"�p�uc�a�<_k�L��N���b�8�E`q�mG�ۙ�d[��=��FxHZ���e@w�.=�/�խx3$EMsN����9�z�P���HA7�S��`�⯅pe-�I�D)�Q�PG"�6�W)��3�н�c|�4�gܕ%���hU}�Ш�<�;�̡_�OE����Hn;�<<-J����%��=g��i�?�����&A	���U�S���y�� �A�Lr�����C��y`{T�(�-�v�d`>��~�s4n����R6���I�Tq�v"��#:G����9�)���ɸ��V$x�ǎ�R�4cXKt�-?��2iU�O̦hh������x���sx��:\]]�p
/��)=<��h9����]D�PJ�Q��2���$#]���t��f��i�q��q���t'���s"�@Z�щwx�8n��{"��CgtkYC�H| �>s!��
�.5�����36N,ŗ��0g��p�����]�Cc����c?�#��d��Q<�SQ	��w��^��JSNjc3�l��1G;�+�P"��(!��۫#�"����f��ݎ���0xOw�pګO�t4�E��f�c2�g���+�9��-��(���!\S��������/���l�F9_����*)�(a��1�����妠�E�q��]#��x�xy��,�1c�2���@B�)'�*T��*�����H�}�5]Z�����\4`#��xãZ�c~� �`�Z�i37J��		/��׽��0��O��qP7��|Ҝ�����!������f0�����ߣ~�;#�(|x,�~�#r�@��b<�t-zOv�L�u;F�d@x�:�mK�{n������C�t�'㈖������h�LOSP��|����6�H��Qh�ȷ0=�1�['����4������'!>�0�����Y� ꌯ�D�ɹ1�Ki��`c8���/t]w�]�~;}�3������d*z��;6?Ƿu�ʫ�꜋���Cp�M��US�����}��*_#�_�SH��S��\��i�dP<��~{�ґʮ���vI8?R+)?��]��3�m�#��yW�V�5D�EU��' L��2���3�ρ?�zc��R#���cS�3*�k寅��t���r��9�B	O����}�G�_:%�Ni�9/���� ��H�J�3/��,��Z��!!�� �Kŵ�Ew���(�����I���߄�5
���D\gd���v����t�:B��?����@�<y�Kh�ʝrR�s�zT��i���"�'���e��f��Z�Y�;��`�3�+n�֨���U�Ѳֻ
wґp�2s���F��7 ���TA6<��C��Dֵ��M���$���K%���`�.dV[9����KO'~������ugR��ƅ���rxT��t�E#��' �#g�%�����87ҩb��zyZWd��mk#�)�>��@�Y�-����[(��O�ʵ�EK���/���_�������_�0�Ҏ���M5u��[q���c׫�d�T��$
�b��Fōt��1�M����\M�Ϋ��p�VA�t�����J����ҍ��~v_�<��D{� �`^H���jR��ԅvx2����ý�L�؋��Lf:@B'`O�Lf e�|
��R*U�ͻB�r�;���S�ʝ�4~Q�����u~3�dZL�i!5��K�Ĝ�������o7�~ʹ��t�?m�)e���m����_\�3�����˞�X�h�1CuFBN��>�
|@眝"h��Ps�T���&_�.i����>s,E�k9�{x�tYr���rO�+�!=~��Y[���*<� �S@�R������4������¨?/�5�ڭ�v��0��p���B��8�p�"�5����o��s�2v:���d��dr	��s4�C���1�� ?d��^�|lT��w�o��������m��<䝞s����|�0�0��1ֱI�y�Cf�n�� Y�k}����>�b��?	�1�p1��sc�˽��o�0��ֵ�ZN�@-����Z�3,��'Z����t4�ǖ�r>]o���p��}�^D�h�ۯ܃�j�˓�eSt��h�Uu	�u�18�&�)���A�3�ц�����S�5��
߮���_�v�Y78�i׽��lys�ޔ�d0�����.�Y�p���H���-'�ǽ=�g���r\��-M��w����-����Zt<=o`��6���=�IW�����qf��Q`��DQU��L6���v%�S��]h��U!�1��t݀S�"y��yE�V���&9�"`<@�.
��%p��xg���U稭��M����P�w-�^�uLc�� ��ARF��i�@�.�N�����9Yr2M�Fs��қ�˿�"�?�ݟb&A�q�L�KP���RE`�"�h?dbT�S�!V���M?�ӳW/;㱝o;����ț�=g��]�`�dލ�
�zl$�����G��|�xܔ �~j��qZS�,nKp�}�=�
�)���GǗG+��q�R}H�'�G��oU�)�ꀒ�1��)m-J�aZ���V+�C��G�R�>�M�^��������`��cQ��iѵ"�4�Ao4߮�B]8�qJa�1��K���t�΂/�Dx=�?��EX�z8�����������#i�pt,���Z򻿭�ᴭ�={��r�d��x=�Cw���R
���?\�ޭE��__�`���S���E�t��+{1����h�O(o:U���ň]�>w�w��Ik��Y�d���]&>��}`�.��C����!�����'�4�L7��S��b]"�Έl��3?z����Й�^dL����"썣-3��l����,6:��xvyL����Uߖ�����/��G�}����ALp8;���T�72Z�x�#T�@���1���A��^K��&Ȅ@ ��L�0��G��p�� �[��F�uQ߶��c佳�)!����̪�幄���k~���s^��B�9�g�k%�_��Ï��9����9T��݁W�g��A���G�u���~⻱��?��	\U�'�.ҞG�0�O9�c���o������T+�0�R�)�A-�x0�mi�7��c'Z(�j����ْ����b&m����a����`�Vq��O��T���tϧ��:�DF�&P�����{�?���"����0�ʊ�.�8��?~礱�3�Cxn�c
�x�ҵ��ϳ>�x	��y`�#���/����Fe��h�Ma�랼����K���
����'�M���j��aM)����/ڨE��d�����h�Rl�{���N�{���ٲ݇A�W��ߏ}����uzt�S�����u�� ��Tk��b^y�
�Ax�)�W>H���=v:�QK���RB]����2��mC�t)�Vd,ċ���O�s$G����[}<i˻��C;���(����?wa�vݕr����Q�~���������@Z�}��ɞ-lΉ�G��jmG�8AE]w�����-F�G�_�~{������#�n�,�I�CuѺɖn��7'ᅷ��{o�O��S�u�t!6��ȁ������Q�����qT���#J��wVJuW��S�v=��i�E��P~N�h��8��I���|#1�Ew�g�L_����-e&��H��6nvy�ZT5�`@����$Lօ�2Ϟ�MO{��N������F�����}s��0�ѫf�p5�i�ď��kq���8����y�.���TZ=	M�0�==�����*��pғ��i�nL�c/V{ ���p�ʝR�!V�����)�BZ0�A7gJ܎EN�`^8T�s�~���h��H�`cy�
�E,!y��>��n|�������LdQF�������P�0&;J�b�r�����M!Dh����jw-k���Y��}�)��c��W"�$��㩥�㹜�Ɓ���_��F0K��/
�t��~�^�@���V{8�-9`�����"���p��W���[y�~���q�0~��J���Ӷօ�cm��ѐ����m����߿x۴���1�ڜd�����^�he�lcq��'IN�׾��2/�5��d+�"�:)뗟�+�usƿxW��-n�����AZW}�y�����r�a��y?�Y���{��iڴ���_kUT6d�f#�����
N!/���Ȱ2�o޵�����`ʝ�DX�xĩ+�c �/�;X����\h+̃���H���\�Ř��1�Z���j��Qwv�g�VZ����	)'�|νd |��	x_�;ǪgoC�4\�Vo��@�7��g�(SY]��"83,9���J+3g��S��c6�z��\�E�z��9���Z���%_��iDf��2�Y�����{���G'���=���x���g:>�;���s�4�M��<����w�O7�p�C\߼����0�Z�_r�[�Y!�9��(���9�5��w�)QM���:�k҉_��e46f�:����d�ȕ.� �.�)�':�%�5�1�{�|��TV=��]<4-*�E���m��]�m��7�=|)�����"/�64"Vt���8sv�aoV��7Vᢖ�]�	�h�>�_�$�/�!����Xy��ԇ"R�9���[�N�N ���sw�%q��c�����',K��)�)<u��ZM�
���t�(گ~�������2n/y}&+���@�y$�J8t�?~X=8��40�sTO���I�Y	5r��LWj��Np�9���^.�gچ�P7xS( Kw����^����=��{����k�JZ)k��OE��Ԋd`�몀�3��}֏��x#��"?a<�0���(��;F��NT�Zd�>�QezЇ_�"�M>�<e�1�Sg1��+x���ķEʓ�-���8������'�`��h^��Ӈ�$�-�N����v8o�d4���f�������1�2�ߢ�{F7v�h����8s�}s���۩��%��׾�Q��f�LǗ�sz�4������[���W�.���M��}�i��Y�a�;��i��=+���.�N���_(S]?�Ӟ��Z�$/
��O""&��w1Ѕ�?���k��6}��q�dx9+�j0�|�ɩk?1]���楣�e�u��P~���*Z��+� � ��w18��u5ie`��]��V�s����$���Ǡ��.�.�p�������`�z���ee)��I}� #�wY��x'+��W�(������&(�{�Ty�7�,�O �\�b>�ի垂%��w�i�|&��Sb�Kz��hq�0"�>`���aZj��Ƌ,d��љL�W�2�<����帪�f8�ioʦ�s�I�gV%�^�\�E�!�|r(���ru��!�8Lf��U��.���'r栍ϡ�?:���v����݃�w n����?��sz;���0e���ʧFՍE�s<�P��O(��2��\c�����~PX���O1�w/���񺾖�����L���V���?����3�q%�!F�<���V���e�!�y���)B��d庌���8��CH��)����9$o���z,��)���$��ft�Y��mlz0)�>A�z����4�{�|��9���ۅ?�ӿ�ڡ ��	�Q@w栝�L	-��{�o���k>���qu��GY�D� ���j��J�Y���<��j�>e0�b��)�q��Ωd�Ob�u�l����s�'>�G��_i��>\��*;o%_u������-����|��B���<ѐ#��D9a崢�7�����2v�x�t2���0�R��g���q�0�u�R'l��U"89�!�5�MB��*��Eٞo-�/(�|�ipǧ�(�n�sH-���#D�巼�*1>�G?X�I�Mo�[�'���vzl��z��kS��� ��o������__����2k�T�I���T���p)X�Rˣ��3��ubA8lzߌ��7�o��v��)s�6Ս0s�»����~��q�w��3��U��OQ���ʯ��1� S+�~-T���G���C��B��������o�)���M����?�Ծ��[�Vߍ��b/ �(q��d�BR�LH�����k+-�WY�uz����Xf-W�=��ٕ�<����;����i����̪L>���BL<���$9����Qm��Gp��:���a�B�+��z��3��RV�갓[��3�gg2L���X�)\�L��1���ǯG$��芦6���,U��HZ�׶j%������	�Ï���r@xc<�S!���@�Nܚ��k��6��Om������/�@�j�EJ�����ӺVp��5d�j;8��o/�d��V\VC�t��S��9�9��"Jpj�B+�[7�K�7 *�e��^�3�3c[,U�_���1��2��z������a8%�~��ş~�ޚ���o��unYr��䶥�R�ؕA*��=����y�3��L���l�n�x8Yʢe�%aC0FD[�"�W� ��!�Y�u�0�q�b�t�'�c^�Ǆ�T��N�i�"�v�C����������C��$�ί�VMx���n�1s4ݟo@'�(2��,��?ZxqZ۬���Vd>�0��u�@Hڠ��aR��U��$� �j������cɨ�^����Xу�S�.��I\t#9�_�:�LZU����a;29�G�����	�ճd���e�ꎆ�d�`�$��g������*��(8���jG�.E��jk	��#�
�L��VBy�S���t�s��H����#l��XU�[�u��m�,瞅Pz�6*D,���.�߻M/NGT�hǴq2X����F�Ά�ﶽGG:�,{V��Nc͜4��5:�GC�1�*��m�l:�z�7�#�\����_���<��\3�Z��<�������S��=<(G��k�0eg��k%Пrn_>�A�>����L�0Q<��z^xa0E*�0���gF"R� \�=ߺ����?g��.��n��S�=�h�=\���C*R��2��p�+�7v2��S�F1b�4���������|ɯ���唻���:�u���#8��2��a)AϪ��Զ9Z�S�D��j��1#�QQ����s|��⃧6G�?��D� ���a�ڜ8�+g�C(��otF�ŧ��4XU�9��X��}Q�����F1��t�:��nTM��{-v��L'J1���~L�*����Y�_32OD?8��H�7&�|�0ٮ!��9K�J���N��\~���)�+�=Yֽ�����<��G����0��/�)�d�`�fh�ԫ�?����N������t�mF���U�p��\OhX��������𻍌~̃�|J5I�gB��7�?B�'�mh��Y���VQ`Թwl�����Mu�ރ�e�B�z���4�������3�M�҉�/Sf��<��Z_���[+>��S��#���h�>
��Wy�����GS7ʃꍻ����WR�st�����<��M��[���)e�/����}-�A4�xs�%�$�h��&��2�p�+�� �)X�R�?g�|��'�,$ZJ�~�p���_�d!Ҝpu�_�a�P��ta2�/�%�3j�/���L~��㗶2=Ѫ��LC�(RKz��.:*�/J�/��Ê�i�ǋh20i=�����`��D,lF7f<J��aȔ��3`xfυ��$'���C7��rD����l��x�c��Q���	Y7|ݻ��Ƹ�Ӿ�y��wɠ��O�%<��7��E�Z�qr)����"�4�H~�amЯ�n�z�/X� ��׼Ə)�߾�w/������QԒ9s�A�`������Y��Q�=�O]�1m�����E��_0��2��8�u`�E.�W>�)���D�n1�~V�R֚}������u��hR7����@!r��͘�6����Ľ����R�����Fk0:�oPT~��w%K�D��0T�"T/=%�c3'w{��$+~=L��&��{��m�3������턒s���Lf�}EQ��lm�2��� П�!~//G�6m��I�����u�4iOO|�[c2ʧb�ǔ8�X7	3��F���+��J���wd�-^*�H<y'o��ŷۓx�]M=�~]ު�%������!N�	������n?J�����^�鋜�Lr���_k��?����mҸ��۠K8a��T�
9��@��5�>w|]�9�=X�cK�s]��?�1n���t�Ɗ�,i�6����1�	���"%����/Eo׋�g����N�ߧt�;/�Oo�.��D�h�����>�9�S Daí��o+t����TH1ָ�?��;��6�|^����A2�3��ެ��1�-��v?[=<_
o9��]+3�S���Cf;Rˁ������bl'��cFU��=_2���&5Y>�)QbnP(琱=[�-�����*j-	�B�I�c� ��x8�G_8�#i�X�U�5«�ZΝ����"��1d<a�S �OO�r�5�>y�9p�z�-QZ0�1������������Ť��������y�h-���U��3�>�r+zE'�\��Ƃgj�y>��� ˸���_c�Q�i/���,Gu�����8�ɼ[��á
8�@T�Q���[�z7`:�W���s�P��Zf���rӷxF��C:�^vu�F�X�2�t�?�1����~�^>�x�WC��,Y�;��ky«�%(A�&.��� ���"�O����paһ���o��?�������\\(�*�/G #,) #�e.�؀�����v
X�����m��D�	!�D%7�m��s�p�RL�ю�<{�V&.���]�"ׅ���(!;� �,k�,���;Bl��ca~9׺O�-S�>�sj��TX��ʻ����]�C�\��S�T�n�Z"��	���K�x~�hT<ߘ@Y4M9֭П��h�B�����U8�7y�{����=r�NJ
���g�8?E8Zb���W�˃W�=h�|ix\����xz8x�C����� �Ƿ	)x�Rtm<��'��Yz�s��XP��d��'�ߢ��U�2��Ѩ��X)�8������ʺ~��9##Of[mt:-������'x���u��ێb�z��c���h�����3؏�K]Vn��V	���9�����O�������`�c��-�/?5�����]�3�
ݱjW�)���s@t��PrQ�v�}gh(�c��������T˾�=�V1x=�T�3�pA�1���P�9&�	bK��oVd�݁��͗�;��ޜ|J��s��9E�"�xP�Ȕ��1�'��k�w������Z@��ȯ�*R9����8�#!ޔh{(�碍��>�� ��׍	��cfj.�Q�#�\���oQ�Ԟ?��~,�{��u��7c��Lf3�`RcV�V���0�����կ�R0ɚ!�~u}��%Ϥ�k�Ms�r$���v���.���::�WJ��������K�֯VG���6(�����K���'�@ 4���˼���MoJx�v6���IwG'�����㢊W�
�:$��DQ�3ɯ+��?nr�9�)>>�ΜA�6hZ}v����o|>����׭Z��h��Ou�{ZC[}1��_��Cr�"���������z��?�{�w�ꏅ�7`V�����$���X՟%�b#�e�{(�{SO)��8Q�l�������y�Z^�E��Ya����u�Dpׯ��{�b���W�����p
����iZ�]rQ������i��vP+�������7��.Gʩ0�w9�QI��f��D%�y��O�p���-����Zp3��b�k|��T��i�Z�{;���Ѿ0���V*UY�O�_&�Ny�&)6�Sǡ_�2sA���)���N�����폽����(C)-��?u~��
i�OxH�S���|�j}Q�q,C���X��|�-�4/��m�*��«��T7=)p�'��_�o�ޠd��p[��[�,���q���҂�k(u!�ڴ ��Y������9�x�U��鶖�xEKfF��$E%�nFt��� �h����@�3�~mL�V4�]Y'��5f�ޛ��l<���J+/P}���#��Z�D�ț�6��W$�O�4��H�����ު����?��u������O��Ϙ�2�c 
@���'7%��gV!�#d�	As�D������*�*&1���	������J]�g����I8��=}�� ��p�@�Z�Ft�����cB�C�ēK���d�ձ1����3�,Q�{�b5ż)�h�w�}������T��� �����2Dխ��X�ƄR~���C�����-Rchd!G�^h�o�z���o�27J��ڦ ���t=�ٓ�8���e����o���U�0#0x�d��u|_s*{Y>�ˣ�A�'Z6��q�oXF���o�pG�}�h:��ѢGo8pBs�C��1�X�j�'�m ;�@?t�%��sQaW��#*����s�Mx��3p�Շ�/��F2����Y�k�ɘ��Ju���}eω�e���+��E@x�48�7��9���>���J�>:����  @ IDAT=���5Y�*�apy4��b��Ӌ����R�����g���-�!D
�s��
`=�_@�S��<#4L���EV+�ٮL,�A�P��&6��T�o}�y�����J�����/����R���Z���f�XU���z=�L@�ǯ��ꛃ#��o2
�1�Q�)N��d8���l���֗�)��S�[O�x�t�Y�E�R
�A9W���{���'�� �N��K�{��=�x8,ge�3Y���m[t�c;������;�+��Hgg���D�F�}3���ف���Y��n�����Ù���h'�V`-�����
�֢��,n���[e�6EN?�ggf�Е�ӿ�炳⡞�}rz1��j#x,[�/���Ы>h��ɺB�����E�Sn�+34Z�׽�V�l��1��kF��x:_�7�C"o��Z��>s4{)v����Gc����/����|�W��GN��[[x�6f0��S��.�s
mBiӌ75SH�Qy_�����i�Wa
����=�N�f���HIg\~�ጴ����eʑq�)�¤ ������6�Ƹ8�Sz8,�^޺{���a�qN:�3?�K U'�Th}��&���b�o���6Ì���q�BĄ�0�0}eZXǧḖ��A00.���'ẃAY�]����~���� ��
I�H���[ U��u]���I��xa?��gz^_�W��ٗ�x���і3����5$��Y�MZ�o�o�g�G�q��Y���,y�}mM�GS�
"�2�?�À��{ߨHI��FE����M��������)�j���#��t&�f��L�7�L�q(3����F��}*u�; �)�����[L.��������4��Y}��=�Lg��:����phl��ɺ�߼������֝��Zs�;�OG��c�h=�$����s�eq��	��ĵ��'�<�1|FO���Ϫ%1�D���綈�}���a��c|a��9��c�yU�sڮ�K�1�����n�_���EA����w���p6e��_����YT��ԉb��ā*ֲn�f,��3?�� )|�y�[����`:�1�����Vg�'���V�u�V�Օ�2��z%U^��b�q<��R\��6M��I�l����>��`<�V�ٺ��˹��9;��(ba�G���V{a��=���^<;gv�� �E����X�w�n�,�Uǹ�'���8�@���z�m�<��.ΎB@?��(��zJl]�n�"=��G�;��Y-��fD�x��*7=e[Wy����߷|��tr����Y���=SƳdOO�!h�z:�+��+X��^�?�����~�X�;��6�d�����)X��k�)B�$��N*�躏Ž).��^e!8�VGN��o����,&B�������F�~-s���S���{���p/�>���
�o�R�p<����^�Bf�q���7z0�>
�ٯ)'��yN�Z-G���=[��J�~ϴ���� ��Ƭ���`�ǫ=����nÿ�G^��L����1�q}��?�����d�ce�W����jK�0p�a�#�����{�U�ǽ͊�p>�����.x����j�?�I8���JV�GU�|�Y!M�Ξ�WY����Σ��3�?}�¬����םL�/«��I.���,/�a�-M�n�J`��4I�t�Bo.OndW�����E
xJO�7>���.�1��j��w��9ݾu�7'ӊ�����3��-���7"n��k�o�2_�]�ll�d�@y��$$&0a����3����2�? ��m��]egUe�3����{#�����#�ʖ0�T����sv������q�J�SA�>錇���Cs-}�e���9DrfG�5d�G��落�ap�����vx��Wp�h�.�=84���^�#����%�
K�����HBAGK��H��lCݽi�>��Wd�<��C�iP� �g[EM2I4@�b�J��$�bH$`G��G�i�������5z�Z.�@[qEt�mM��U�\ū( �E\�9� ������R�C�@�ɯ�U�Df���5Exh)SYD�%���+�<�\��`E��O �Ko��h��G�5�
�e"��U�xM�R�[�U
_%�EY}�n�Ì�π��:t��M�t�,�_xH�T-V"�q�x�t��gK��2i����ҥ�0Bn�U},#�p�VE����gh�K�w�y��tqwp���C&��^v�
k�$A��>Pqv���ۤ2c*Y)Y��
6���jJءHT���yl�ᅸ���Z^IA�U'e��jO �Β���t�I
�c =�G���������~��-��W��=b���XM2�`z.42��`�zի�T8�V�T�sA=(�ė
�u	#�~w��y�UD,����Y��j���Q�2�U�/�ٻ+y�Pԑ�6�RY���%�P9��x��c`�q�v�� ⛱�&J]5@Uf��7k-�E \����q���!���gi�-ĺd�P���.�Ɛ�8H�47X%�*�$��1��U����y֓u�J��^�)q&��\x�A(�Ma����1�m�g������gj�kt�C3��E$���tѐٖ�|�_�i)#�Ck��&8�Y�&�"��,�8�L�-gH�h�Q��_�9�e3r��ؕ�+2�E�8�� Py�)x�����,��aH�L�k8 B�ʝ��^���e����u*&7�բ4�F�1ly�1=un��*���F�鞨�E{շС��~��.���tO5̅����e�{��b-��s��$��6;eXZ-_`�t�"�I7<n9�1�y�!Ÿj.�BC��?��\.��r��  .�eE�}�D���[�D����אG��*d
MA�R���1&��d����-�y�bP���| �8����:J��^Aap�n��Cq���U��� "o&��?��6&�-���7�~��P\�հ
G�^0o�2�ʪ�JJ`��K-���*e��_RB<)0D��
�Co�T���ԥ����zB�n�lO*�[�^Zq����ƞ%�Q��c�|NRí��YxMZ�? �f��M�$�,��h (��:9!^!�W�-����w9 �u�l�pBҁ�����5{�#�ZA������<�B`��҄���)�e[՟8%�����#Fg������x)4��H<�9|d^�q�vD�Y��*���@N~�rml�Ӯ����9��;�v�s6ӹ`,;�iHy�>g����Z��5n$�S����/[a���e�Xx2mG�r��L�S�DQi��xk̜���P��۩��~�),*-5y�F��*J4�a��C��b�dHp���#܄)�]z1`I���H�DpPD0�%��&�EPt�dF	�y(K΄]�NY�%z��g�q�널d��� �F֫�F��.��`�)��x�W�Yg���aH2���g~�|Ǣ�
��Iyz�$=�[�� ��+8�k��Q���[ެu�f��Yj�o�Ղ (���Ԛ�G��(T<.��4~�V�ض?s*F�NE��|)S�.5.�i)���:�	�!̤^wzXqzjϋ8aє�͔I{Uν%��7��S#�UN�" ꏗ��i�)-�sG�]�;CA�����^lt�/�t����b
�*:�*�18]"G���]�s�o_�2�3T�3s�䅢��:UCa�C���ܧ���12G+?��ZY�B�N�A��S��0�PC;�S�����B��|\����7>P�q5b�Sck��z�٥\�9���~���"a*:�
n\m� 	"d|��fF��Qw\ӕ0S�H��T>��.[-�|Q���(>�Y�R��g�.��ƣ{�շ�O�)���+e� p��*�a$.p�	�.)�iTJiȗ�\������}1�X��$gR�
���T��F]� ��[�������V]wQQ~�
��F��Ɏƶ�����]T��j+����#���}�t0n������f8��U�zP6�q��V�B:�օ��
d7m����`��I%V� �RG�w�2�3�ˠ޴U�H;b�#�>�Ve��:1�)5U�K�zG)���09����5`�c�Lֹ��Tz�/�����ו�%��2���v�e B�ezb���8�� {Mx���o�oG.J��A%��\��T�I6]��$�o�.^\G����q�ދӛݔ 'U��"a�U�ԅ!',�.�O^LH]�س�4{�z1��C� ��KK!~�#3������O1=���> g�&�l���ߌG�֫"�cW>x��u�l&�����(Lm8h�4�K�n���,�K�)Ѝ����5C���0�Ϭ�f�[�T�kX������C����Ѣm�U���4�y�S,�ֈEy����<PG�3�憻WCpѠ��Ju �U��Ԕ�qX����3B8��;��=�t*�K�#�VʠH�%�<�/,F�ţ�쵝e��w��
��w蘍|��Sg[��ȻpJ;�I�ŝ�He� �|�k��I��"h��z��m[��Az|dT�Ĳ�Lz�9E�('l����ߴ�A�-��A�r��,[�@0'ɧ1$W���;�P���#���1�[;�����]h��i"�#�ku�h�h\�oc~�|���0�7F�]���M�~)���c���rZ�p�1�Y�F���/0*2$�H"(�"K���6��PE&�JT<ed� �0��R�b�\��:��)�ZDR/���:-��*�u�G���E�A�9�>��&Ƙ�]`�drO��߀p�=�F=�����<�[����^�J�1eJ���T�R���3��T>���W���V��7$��O1e�N~I_���c���}��3�ʐUe�N�Pe��iL
���l�����<����`��&�y9B�Y`�g��v~D�JGY��<�:87m2�qy׉��CDa>;?��ǀ�!��A2U���U^A���|IG�m���ю�-�qV�Ǹ�TH�b ���a��3� ���=���b�ve�<����ܗ������I��N�Sy��G�i0^b7�c���=�y��?��u���2�[���($����� �s
�;=`,��L'�o�ʉL�FY6�%*�.��Y��^$���(��7"x2g�a����A
�k'�c+��ќ��I��1`z�y.��5�{�O�*���U��m�zJ���B�9}�h1�������I\5��s����^�6h�6s��h'3C���W%,%̅�M�4�=�xRG��n��ߺ]��ٛ�=q��p_r���n�3�:��ab��U��W\b��[�(c�3�J[vy�zyc"φ�h���v�\���LB�#�=X�C?�TN#�^-P::5I[&��JQ)�uV>eJ��Q��G�<S�z xȀ��o�	P�4j�W�M�Ugh]*w���Þ���`w���Q)�Efu
�=S�~�#�	�F�a��)?�\�Tz*�Ze�1O'��>�֥?�.8�@뾾�m1��o�<R��\we�2E0h@�\�ĝ�4�v�|N=��g�
�P���h�:<����8���oY���m�6�d�#b��� �eG#��cd��T��
�8�?�f=�"���ɞy]��v<h@(^���k�J�0���r�|��9��~>���^����܎��m����(�I�����J�mpu�u����1���H��م���F��|��t�7�VI����Bn��6��G��YYH��g�#�A�(z
��XB�G]O���8��
�P٩>�>5����`{ª�4ho��v�3��k�Y��c��S�c��Hi��K�2R*��<. ��Q��*Q�^m)��/C�DIY�yu"t�)�U��Rm����L��_�ISڬ��"��O�$<!�?���E�0���
���W�Gנ�4mi�h�:��;��
.\Oİq�VYs��E9��-�4���� "�V����If�2��Q �T`�:�}�KY��&#5[7��ڑ�Z^�nX�0� Ҝ���d`=9eD��Wr����aM9��ߌL@�s�����!��#��^@
UO� �����t*�(坱����Ѓ<u2�P��C����f�dn�C��2<1@,�d��x�q0�
�i����5L*
j�c	(x;/����֊64����7W�#_�	��ܑ� ����\�ц�����P�k�91hl�����$����MY{|�.}h����
�����8�#����X�i�zzF�50������!g5c��k-K�f�y�*���Cӊ�A`�}Y4��ۙ��-�����h� �]xKg��	�Ԁ�J'��kH0��5~ҡ{ �G�D�@���%��oӮ�S:��1�TA9�;�(�i:�B�$a4ؖ$�G�}��q����#
���G9C 	�{¥e�IFRVA���c�q{=EֺUᓁ>{U���� (ԗ�r0A"�Wa��>���q�,O� Q�/o0�@.Йyt?$�+0�Š@��{7�Ḗ譊ާ� �_VBN�\8;�:(�̻F=3���.��g��^º,o`K:)T�.	f2<��8��)�.�N�ÎCe>�ak�S��$�4z^��Yq��BL���"������ ���amD�O!JO�ӜB"����/�P�#0E�Sx=������njDp�!U^�C�
~z/0I'�YgAu�'`�_
����f�(偐l�`�"򥋒3G�Ie�������'�4�*�x�
� !m.-�{�d��|�0���q��W�r�(�F�!�Lf(<���O�a��3�r�b�c���4���+7ɠv�.�ll ܘ�ϳsegXD��l����AZ-�r�iM�$g*6��ux��Cc�}�E �U�V}�::�5��3�*��/ZU�X�wx���W�̂�@�`/�T��<w�;�VO�!C<(�X֏L��ah#���M���hrq�@@t-��zC�����9��cܧlۥ�0�}�Q
{B����ͮa�եF>�^% ���G����u�Y���~qy��ӣH�߮*te�Ȁ Qr��s�\XVy��o��d՞��,�AJ�n'9+D�_o�ʠi0�>�ߔ��!��]"�<�Ѻ�2�G�J��!�ڏF-|� ŕ��|	��	���V��Oԟ���{��A�z.�Ҽhe7dg�j�h�����q��� g��=�8q�Y ��>�L��#�vL��.Jօpr��u;K����P'�As亼ea�^D0ڮJU�j�E��|�Q6�\�
*>�ئ�w�jc֍ �z9�@ D��l������"�숏�����J覜����"?���cɪ��>�x�+<ʕ����^V<v�����ն���Zs�[e$4����_V&n�Ӓr�O�2�Vv"�Z�гd�n�/�Ho͕�+���I�c޸�}�ʝ�i�0 ��G�tSP|hD���PF_W�<5� m��#)uLxҮ�5�C|6(`1�ZΖu�Ǹ��#���pL\� ����uM �wrF�"ӏ6*Ma���GLa�u۳Q�+G%>��#���<��8I�����r�T���{�-����Z�@�pu��>�K�^��{?�}�v���40{��a
���y�>��4�v�n񪠇�����^�u*�dEm�Ŋ[�c�#XP��ס�<�<xG�!H�	/"s�m��w��ȣ۲��{�� �е�:��7I�tPT��ȷ��P.Py�O �K�>|J���\�萤�2�)�� �L��D�n�[D!�XKM���Ax�g�}S�ir�K��^�Cg5�^���.p�D��^G�����v�un�i�F��zz�%�B���e�Nm++�[QfG�T��@��P��B��At�s�m�&p��
Ep��5���"�HBq�o��H��v�ڦ2�CpoI�P[-����4�{&dL��V��������
�0��T���X�*�!��o{�ץ�T"=�_Fz��m#�j��0{���띩��?�C{a��fH�O���9���*��+���Y3�!��盔5 �:�L/F_6<���U�NN.�=��l��E4�����LhÏ��g>��֝� ����kzY���ӛq�u�)�P�@t�S7n�R�'�L�ߡ����������'�BlT�JA�֦.�9�ŵ�~,ѐjҎ^�Q6�d�u��LLE��L]���[;�r�;[�C/T�l����lz���q[�XM�boӿ�^�!d���wdHa���zτK�ˇ��g��[�F�p��)�Z�7��*	����%*b��L� T� ����%�U\)��ZKc�<c`2�!�[f�-�0%I�=�v���Ѥq�d]��8x~t�I����4���>M��(eB�m��$9�0�1n\N�}򒇊�-d�kf/�F�K7(�x�WASp�R��̛�� �z�Ps
/��\�v�z�f~�o��#�^ޣ��=�'oz�B�K������ph�(�Ճ0�ty���ݐ���7g�{_|V���pS��c%A\ȯ�"��9��߶%��#C� ��:�Le5��D ���dM�/x�_��0t�ٽ�Z�m{zS1Kd��b�ci[�����������7�䳉�n��L��N�)���	��|�E��<al�`
�=��	gɞq(�.���:u<���*O�M%�g���uo Vs��t�ãUVV��A�ϝ���ue���� ��Ҧc�M"�QF�T�bD��0��� �i�"��L���=�1
]���[��^�@����Ȭ_0@�����l��N��M2�]��[��^G���� # "�n߂��V��F)�0�TͣKOC9�UC
�n��	�Uɾpp��L�"2$�;�sW܄�ڌ�(|�#Nu�,�3��8�'�w1�|�_�D)
�5*��W��2����^5,�2	���͡e�N�5y�2Z�s�⬰�ҖȒ�絸T���y"��)\�t<���y���\�SV� ��x^�\zI��<���R�t/)�Bv
��ˠ�2�1�cg��X/&Ń_oS��@h� π*| �Ǣ��/mas��.��cD���S`�|F�����&O�ˀo�����@�Aa��u�����rM�=�_W7�"�	Ej]2��a��(�E��NΣ4��f1��aL��T�UF4�6aO�2 +���G����W���]QV�aDX��o�r���T���g��v��r,=�D�b4��b���^ø��{Z�nZީH���l�4gyc
�uG�Tf��S.V�k{H�őN2���^���!�Z���/��k� ɦuA�\x�|(+|Z�d�*!���P{�P	K�S�1�$�~��g���dz�(����%#�X�N(!��t顃��Zr�St"d�h����T�(���������NGVh���f�>0,�Lmz��+AG3�+_9M[^�f���0��5znIȗ�@啿��0h�'y\Q�|ӓ��l���;�C�[Re��&�0s�)���]���;&<�j�@�)d�-��GR��i��#���V7�m��1&Ș�����	%W�̸ŵ�O��	z��A�	Ϲ�1B�s�|9e/�	�ڐS�Ǹ-w�p~*P���d� 
�h�z�D�)� ��=|E��7^JOa�Y��Q�ܵ? H�h��'��,a��L"�Z�8���q��jE�G��ō�E�]�L��&�Nq:��8��UP-8��̚�0�n��'P	���!dr���\�Iöcd����Y�5�)�塶���a�L���D�n���JQ���>�z�나��HS�����ĵ�!hy�R��6�x���vlТ�	�3�/�w����2��Q�x�m�a,�EhKasX���2%B��@{j��0S]`�G�<�i[ّd��i����>׫��
|��e �^����@�R��yy�k4VS���u���pٛz���+2����dhb�m�.wů�>��ag�:��o�'��N-���đP]]_�5��޲�|�z��qi�Sh�m�n{��/��#��'�,���Ef��̚W��]��qbE�P{h���D{J�K0l�gԟ�L*��hQ�<��}�
`���XwL�J��*��*d��_���� wx�-�i۠�HFBt�ղ�Gww/���\���e�[PIzP��
Ahk<elg�I�d��!@�����W�g�}����00u���N�NT�/a�n���S-&C�]@L�"&T0���1Q^(Q"/�e�\oP��o�C ×!�^hM�֧j�(7�Je�U�$X�M�f=��1Z�hU	����F�h 	m��hFEz9�G�&v�1!�h� ��yʊC��c��s(��YsQ��ְ:T����GnA���ͳ�h*VT�[B���)���ԧA��B�� nm��"'�CG)��%�I�ʘ�I_"%��+?����8Ov�ʠ�Ӑ1�t>�[|l?�H�"'�QG��ʕ|ƋG�2�pT��(8'�I�u�s:�K�!�W���S��:�}
�eM]5@W/ɞ ������ۗ簜�
�U�b�Z3�y���L�_zBn�L_��H���ވ��}� F�u�b<$&e=��� 
=8 k��f�AM��gE���r�������ʻ,����J���t��G&�~���7�2�2�I43E����ˇ5(�me�"��S�XZ2��1tE����w��%^�=P�Xf+�L��I+SyԪPS��6�)g�S0����18�U�� _ա�)8��Y&л�����A�@ �3A��=f	�=#8Pq�aXh泳(��Y\�C�2���"���H��%��t0(R�W�9A�YFeu����Ѕz���HdV�s ��T> ���[E�ogM��<1�ͼfW����ܫxO�&����S����������O��b�v���)�.�a�F�xrD9l�u��g�!>t&�#tRoi�H+����M:����%҂Bu*OlF�oI*SuTp�]�;�\]Xd��
�&��^�xx�R�:\��TUB�Iy�/E�W��n`{N�d�!r�]�rsbZ��6���?����b:��Y QV�8�XdV�p��_���W���p�;�[S�*!��Np���
hq�(HQ`��T�&�$�p�W��v��4.��]�*K�K�4 ������M%��`!lU���&IVg@@mˑ�#e{�in�R0����'ͅ�	�O��ZL/�e��[�����=�����H�и�u�nh%O���H���sR��+����Q���,�)�d��m��B�oȯ@
+������FiNy��>��E���e�W(�$���˰�B�Jj]$�2���(J#m��^I�Au,��?�b��%�q��;�*mV�Y5ӆ>�j8�����J�L�!z��1S��/0o��æMnZ�4��J#蒊f��V��q5
��<��)�±�r�E�R@�x��@t r
�\�H�â�Qhdr��3\2�̲W	���^Q��a�S��0� v��QQ���K2܀��P�Nz��`��a�A-�h��A������Þ%��]�^�]`(�a�!����Q�ok�(w�p-/�U]Y��ǋ�=�j(�k�9����9�0
��\�씉NR�yK����s��6������g�9� �ߔ�cy�w��hb`bS͔���v�/�J�,kN�g��p�G�!L*H�ɧG�����~� �")�z
���������2�.:a�P�S�Y��P�sA�G�$�Ʈ�Y͵���Gi_2T��q�U��C!�SFyfW�y` ]ކo�?E�'�@}g���65�£�����D��J1�L�m��a?kUJP@Y���
}�=BO{Ki�T�" Z$ \c�^q�^{]�L�PB��q��U�����Kd����6����XcǶc,�ʹ�da��>� �H�o��������3�0�ŧ��U� X""�sn W�t��	���E74�C����a��������&.Ρ��S�6P���q�SQun�s�BC�Crǿi	O��9$�ok��=�ϥ���?�h� �*���>�(��ȁ�h�����.P�:mY!��5�T/����˪=KqϏ��}*������p�T�q�2��id��w��Ye�DU�ݭCO�7N��E�|�9�r����N����qJ�ˋ����~���Ny�xȂ� y>�-u�oRn�[F���Д
���D���>սtdE����w`��(�L0D��/2��0yV���&����UX���՚��ӵ�ɶ,3bџ��B�1gBh5��K�{2%��9��E]p]᳜��.�����MF��w��L�D����FnK -:�\������	SHY�H1$��7<������A:��X�|��W�o�%��fl	cIK2AE�B`Y>)���E�p�p�.�H&��QcW��nz
��� �V,cL+��UG�ax�s`��ش�^�+� Tj�?��Uk�_��I����r)AEib=�d��6�C�J�R!l��n��o��o[�3�|��6�V�ox��2�禂1�4�yy3��_y�X
�����G�J+�m�B�b��K:!���R e�
��?K��a!�(nQJ��.�8t*����}�4�

 w+]95L��(�P2�l��� 4��^����@��e>y.���W����(%��MR��	.�e:Щ���5�'oģd��Y��>��E'��O�L�G�-�2���g��S	t%��˾	��*x(�#+��:`�R�(�-�`���X�,[����$���_�=�an(ɂ!sS����B�;�:�y^�x}h�z���%jC%P�"Q5fQ�����{���nA3��Ş�l*���[~�AT�
��v�+T^�%���V���R��	q㗅y��\AD�Th�����`lD�H8z_�[^�t��e�9�xM��ېJ=ɏ ×���$�4�Y�]�e=3���X�V;e (��rMp�aƘ¯�Q�Vrb-*_ ��q�*xn'X�cޡ��S�@9=U�����Kt,ưh��$�ŅV��5���|հ���P(%AC����BۑK`���G�jP��e��H�Ju�R�R��n�#��:�4�H����	^�-�nK�T'�.��Vx8�tb����`�&s����).?'���]PF�8ղ�h�u@/�g'Υמ{w2��ux2*�ӑ�����媞�P��dz�2�Ld��
�v��`)��#���`����/=�A��$*�m�a~ga��]�^�q{��,�F�|���
�L��䳎�ؾ��.���.$���]���*����Ƽ�L����2�f�C>X.u��H{*��fH�~-��szb������5�nb�h��&9N�1ډQ�y]k`���Ѐ��b!�-4H�4^�����E��tq�}�?�4��za�P��}Y�|	�H�рo���%��A�6��p0��$k��s��+�������}=�R��Z��R:h�AM7�Ǟ��fG<-ԕ�d��,��P�ɹ���GSk�FN4��U	��<��iCx3�Q���q�:��v�	����mck��mnQ�S�R�-+���P�=1ɱ�$�[׻�@H*��ly���Q� ڂ��c�Y�~��\[�X$���w��N�k�G�����D4�(��/F�{�%p%=˻���:[u]<�z����d\`*x�7��
�	�P��j֟�Sx������\F��Sp	wր��C���!��o��r6R3�U�u��0�E[˼Cq�I��xSp:��3x�ɯ��	�������:Ç�$4�:06�NOy��W^"|FƢ��O�
.%+F!�UM�V�(��ǌ��˓��v�G�P�u ��z��}?qO�R���PW�I+r떻��3\�e[Y���^GE�n��$�5V�"g��O`���-T�|$���*)�����G�d�/�h֝�D�h>�X !U>�N�_��߳���Ovk��H��`�(�zU�B܂���H8m�����-o�^��*�n��@�epbM�8k2f`7�o/�r��|LO:�H0`t�f0RA�n�g�b�t�xH��A�q��`<���A^�8���H���Z�@Y��-,º#��`�7�R`gؤХmHT�}�ɩ�2�:��m��݌��t�S���$16���F]� ��EyV�w#�ƌ���!fp*��7V��b���(<46�j!��U�$�0eN�������B���tdX��Z�:K{U�TF5?C�+e��-h��0�����Zζj� ��-H��v�C;� �e3ʆ���ꥑ�S�<�ļ�4����-�P�2WƓ�.�Gbp
,�\���)��S2#+@�AQ���oh�.�RN���!���M�
�����:�;�{!4������5�Y�t-K��!u	4%�Y��?y�	2T�Dԯ�C;G
���	T�at��>��Ս��ΰ�u�7�	��5��p 60@��)|�4�+�bfi�+��i(�.כ�ɪ�6��D�zK����.��M�k`M���%�i R(x��Jxhe>�W��O�]/¨v	_JP���
f�'.$����)�����SJTǓ�3��N��U�8S3M
Q���El�s�.>c�"��T�#��|]��<*O��pc��ÃQ�V�;�6
?5I��S����L1���R�И4��FJ%�hUpU�R���pI~r?Y��ȱ��G�A�� �	��߻~�4�G�4��"�1�~��4���C����������cr�����Xvq.Z�Iq�#(ٵ�Nh�ը�C6hF9�%�KN%�] �i/2N���c4�]�}g��3p �W�@�5^^�Vy�^�uJ��d`O�濝����$ >=:�i�K.����X��	�JE�,?��]/���}Τ\��A1�6�S�f�X+�jr&A�D�iR��P��Y�%�P(�eu��@�m��,9-�|�>�I*�/��Z��� q'2Oh*���D����P؋��⎺fa���P-s���~]J ��k�c\�	�5�)Gr�,�SAĪ��(���d/	����0m��i<T~�3��神",w�C�wC�\[��ޑ0GTxp��b<t��<t�#��p�+\V���l �'�S��J!,��b��[i�b�N��Y�kY��(��'W��e���H5��^���]^�$h-r�2�����]��9��uX��i�TvBS1+�c޹���>%0�s�l��r���A
Ե�5N!O��J��x����6�1Բ~�%/����7(��8��0f]
|2u�|�r�t3!�#'�YƧsN~"kT��'<>@��bڌQu�a��h��~0���u�'`���3�6Hc^KS����W_)h�>��qg��l9+~ ���(Ϻ�^s��D�+��[�څ���p��/a�I8>l("�u��GEs�����!��yb4>f��������2�Ʌ?�����ŋ[��QLW��Υ��(2J$|�>QRڪ!E�l�О4�3 pƉ	��y�Tf
���J���5����<�I��rO�4��4�g��y#Q,��F<�'���*czEJ�>�ң'��)�Ğ>[��I�^����
�q��=��������;;>�lU^�u��}pn��a��nJy}�
��C���P��]�/��,�!m��1}��i�x�ƩwL� @�֓+(��Q���̬h���@�<$Lye!�8-��4e9 ߝ����Z=��N_�p���A�����#���T\��A�c6��p��VV��'J���>H�zc��JSiR �Y�-$�!�s�d-�H��� ]��2��" �y��]�B � /�4���+�T!��H8@�АEx\V�|Qr��Ek�L�n�n��W�zӋ! � <��O�B�<	N��fvC�"U~i��І4�y�D%T��c�{�aN���L�a��@���nE�q��꽱�@���W�3�J�[��(��&�[�H�IA�Ŷ7��;����a�ھ�J�\G�{~�ڃۺIA=�2ո:?�ۨ+�)(d�71��z��
e&�Ҫ(��
{��i���Czp�56vB&i��Y\��hX��Mʧ2�8   @ IDAT��q�Dŏ��S�pF��m=^���H���:[��y�<��&D�[
MWD~hn[f�o=-�U'>`�7Ovr^a$:��mT���q:n�<(|���w�H����ܓ��_u"v)n_�_"P�7���"o �ȹ�5VN��s�`'�5�*�=DrzΔE5d���D
�LQU�"B3Vȸ\�K�����S���l|�e�Z�-�K�Tg����;Q��&ȩ���I�yɃ�)�5�e��^V��W�
��u�^�Jhw	������J�ށ������b���A�9T��>��^N*d��:��(��1��8�o���م�&�nس�HX& ����V䣾��i�?~��Q �B��qw��t�K�d��Bs�]��w�(�nL
�(�3��c��Krj�K��4n���>�Kzc<>g�=������4�n�7�b����K���E$2��`,�g���䤂��p�sh�2�q���m�d#��W�f�&zⲁ�f�n`���@�Іڇ�3�ܑ`�y$�F�&)zH~��O�z?���l�y�G���!��i'��w������4V!��=��G�"Uo0��邈��2
b���.�ӛGp���(6�8m$l�P/@1MJ6{�bԋV42_\
b>���hH.׵7���+ƣ(U?3_jԝS`��&��a�� ����}:�&�#�9+���z��H#�����PS��(9�"�ـ��Y��>s�WmS��r���A��zk����l�\��.�&h��si��P�t}��65f�(����@��c\yC0�&��*�Y>8D��%E�?�G^��&$A�>�乒I�-*�\ �j��1l+O�|(�'�␂g]{�7�aP�s���o)MyWJAh�z"_�R^�#桻S�˳�NQ���x[���1�q�����Û��7�e�i���H�WC8�!�_i$�E#�uC]�L�=�*~)����#��z��޹�����)���e;>b�سW68�ZH�K/G?3b�F����QN�%)�2#�a D	Rgy.�\7P��
�P���	ܡ����r�7[)�-Ä�g�7��z$��g �Vv*f�+�*k�Ny���F���]�`�&eK���˾�бl�aPItq���+������kK�l��V���ϡNzg���rpr��J[�>�z݋rG]I�ig������hl����h�R�Oy7GO1��'X���&��Kh:3��B΋ey�e�ț(,e�[V����%�րz};!!:�,<�Ӽn��F�0$U���q�
;Eq]����1Wj(!W�*� �a/�)�ѡ��9�������1h�Y�JX��D#tN� �'��������)��ķ�Wb�
^��U�ӣ�P�;ﹺT�E׳b�T�fܥ�w���ӎHx��=?�6�8�D�R*x�2e�&e�5DƸaخ�2����{"����c�T�A,����3�A���� ��9�EN���6�&�ThO�a^�U~�-nP����?�8��,Q	��zm�8A�s��
?��B�H6���,�0Z �!�?�)��U���mQX�^���]���L����.r��&�UiM�oN6�fŶx��r�+."r>��"�e`����Va��?�^�0y�$��O~皲��Z�Ǉ��z�z��WF��d*8�"�D28W|���jY��e���GI� s���?�	������p5��83�@R�=�3
�|�`f��c=��)��b!�; ��:�4
��5j',4KOoR�CV�id~ň�Q��3)!��7q�cv���{�둎T����K`��#�`����J0H'��'u�?FzW'C������k��V��Zʉ�Ň�%+�+^�W~Eo��:#w$��2＆���Л6V����af9&[�R�!�rE�<ۑ:%\5]��t@=���Ci-_�J�	ؔ� ��=댐G$�BW5�-E�<��X��*���Q^:��e5����L�+�,�����?����	�����CR�<��:���:�h�g����,3�X�1eW����(!�Yhت'���}�25J��Ld��x>C���h5�H`M�t3�P=e�ŭ���I�W��Þ����rSO��y�y������Az���Ny�s�y���è�)Y�$n��<��zW�A/��P�Ó�K��������(=�!Q�A��q�k��0S�vD9äQ�Du���s�m�)�t|���e�j�=Jo���N�����R���4��y�K�P@ĝGᕿ̠�r�<5��������ՙtZς���`O(���h��AfP<p%���>$F5�7�
����b)��+��x�J�;D I{�"�����̊!��H2�ΗU�3�`.�P�P/$/9I9�j�DN�%2y�s�~����%<��I?ԥv���\y��u3,J^`R�jh�O���X7�H����@�{7F n��P�o��Dە��I����1u+}��,����ScQ��JZ�bf�����}C�Z�dn�p*x��Z�U�A����`;*�l�v�C,��8�B��g���LeP&�$\���1#y,\Ḹz��(����|���߶�w<�"��Ku�u-�(ďl�ap�76agDʫ���nc�#��BOD���t�D�m��cl�G=�Sn:-��(>"Z^�κ��A^���JJjYaF�	��0z�M�g�Q>ц)S��<��z���	}��pM�]ɾUn������;QaQ��;�	�8�ӕ���cH�eh�j+�4�vI\����'
��0��V5����k�w�G\d�M�@�e�pcc@��rr:H�2�Ie�P�6�~���@)�^�35;w���<	.j����SX"�(��̗�p�x��pƠ�;��^�{*���n�N2�B񞄡�w�U��0�G����P^<�Hw�e�X��FKU��[� -�~�&6�yU-��ڿ	�z-�d�}���
�u[N���J���V|���z�`[9+�-@*��WR�K�}�� ���۽
���� ywf`�:u�=p6��}W��4&�@4�(��	�4��<k\��Y��ye� �t�S�rn
+Ց),����ܳCݱ�%�U�W*�qJ;=2|�#�P**9�<"�Ay���<�NR/�h-zǭ�D��6e��_T����X�x��U�hs���ӷ��T�p��2���x:��ʌќۄI*�^9�������D��P������K+J�ZϞ^c�o�I�,�����/��2�:DT��M=�f�xZ�W]Y��
���)<�A~E��&]Uh�$.��=�sVg]^]p�f�)%0�^��/��f0�r�W�+BOT^����;uEۼ���u��	|�_0Z?�Pv0r@��28�]~sI{	Zy��Ђ'
��G٩�&��C��<�@�3���ܳ礑T��{]S�~�;:�5p���6�W�X�)JbE�-�b�l����'�Q���M�Gz�|Cw�ҡVhJfq�mgx�v�>�-�]Aj�Ύ��UVg2��B+�*�퀣��a��ո3��'����h4j�Zt��y�&���5�ך�F" J7`�s�{�ͧ��/_����lhl��U�_^k�B 0��N�xY�	�Y�I2�I ��~��͠��1Yk(��͇`�aͿ�0b�HB�Q|�����3�Y�Z�`C���j���R��2;�ʭ��1%0����`'X�(Z:J:�^�L2ݔ&,�i�5o¯��|p�Q�X�$ʋ�/����c�2�Ac~bT�'#K������e�}�u��I��Ǉ�Q}��"!�n�)�-B<K�D��c��Z=�*Y-��J�J�$��ƥOS�h��5�?Z@X�'i ]���\w��Sh��"�v���,� ��<�p{3��T��~���P���I��Q?�zX�������*� �<���?^Q`�𸰮{��r��75FiT*/i�M	�eL�c��Z��s=Q�$VimJ����+c+2�������5�N��}��>x�3�k����׼��
��$���&w%h��z�$=��>���*5܃qY�@{�Dh*�;���9��}�Y�s��o��%z����BbJ9�)"X�oS1���r�Y��Z\�>�e�.a
����(�յ����wX	']Ud��Y�'�������	2��)(�B~�c�Փ�R�^� ��2o��5�-����3i"||(��s	��N�����9�GXCS�"<%|
�e+0���+��G=V�ّa��O��<ޗ�	gM�eև �/sN��w��|=�靡U`�F��N<�� ���g�}ZM�*�ls@R��c�r?��z��m�Ut)|<�4à��w}��T4TS�5��kt<W"��|��h��[)Zz�gz(��b��J]��m�2 k�B|��|Kz=� ��`���3���5k�q ������`���Tu)Y�<g��ka�IY(���������/7o�Qfe/e�]�0� �����N<;�k�;m����|���u�~�Ic�ȼ�z��r���&�+טWB�B�̰�w�����Pl(���*�R�z�'�k��'H|��oˈp\;��
F%D��7���`�b�aP�0�
ƍTp��?���@�öG�������m�'F�E+�ε.BZ���JGY������,"`��Θ���Gߙ�����ҿ������U���t�3��\�]�eMq��f��cu�Ɯ�x�'��Ϛ������ME��H>�l�m�.���ܳS ��d� ~���<���Xyj^]7lr�P��pa�瀿��o��5q�tQ��
@���� ����6��)t)z
���N���3�&�K��bM��ۥߔ*W�	� g��<RQZGNhǩY�#e��h%�䧗����zM�)^R:�\�;�_=[3A3��(�ƶ4���{�
3�%k7n���]��{�]۞��.�?��I�o���1kM�h�ѧ�/�տ��^����&���h�ղ��$�k!�*s��t��Q�Bd�F#��\�W�P�h��D.��|��6u�,GF��7Q�Dʣt�̴gN��C���b�=It*�6�~�o��9�
F]����U'�՘ #1�_�"�v��-��=����\^�M���|,/����
)�Q4�/���|�����,j���\�8�q��C��c#���P^e�&3QҺ�HoVE6�?�%%'�&��|�A�IE��Z��D}�+���7)3�;�wey�N7~���{ʎ��'�����± ���{Q�<��Ci4z����W�W_�|D_HO�}���?���p�AV��X1�g�p��^gA��t-/��I-nuC9�6��\���\���'eMZJc?C�:z��'�xη�ʌm-XR�<�Xɷw��	��I�U��Y�����M���훿�u(DT~~r�-m��ы��@p��P�3	�g+�P;��1�^�ȏX���%{�r��Z���F�C���5iI<����19���@5H���fKP�]���g]/߃�[�-f�q5c�H�D���D�Qƞ�ӥ��P(���uf������*��BcK1�*������%���!�m���V^
�2x���`n��ja�"��1C��6���9֏o�!d^DK#����@c��@c~yc*��OSUoGa���=|�F�3��I�m$��7�LV������a���AU��x\i����$CS7Yd�7��|����t3 8�R�;� 3^ң�(���s%-2]K�cz�t(�sfITM����t?C�������hOO,)PP�g�NuC��$�_'ڑ��(]r����$�i�1�riP������a��<P���%�0���o��G������j���I�z��m����+��6k�v�W'l�<�? �}^)�;����"  6��G~+h(�I����I}���_��ƫ�e� �f;��r������V��AW��2"慸���\�<,rT��q��Fm�k�U����0����5�N^_� 
���n��d�x$��ߤړ��,��⤛L&;hO���K��Hq�ҥ���?У��CN�
|F���ՇgWS|գ��g�J�F^\3�@�ڪ|�
�!�E�R9@�*�a�����1�7Эh�Ǒ�h�m�'��g�_�Y:�����Y�9h&��#,i�!�Jn�������o��d-G����	��y���g���r�����x�M
���"���@o#Zo%��rY�6�V��E!�=�N��3��	��s��������$�!�9��=t����Ȅ�R��2��2�{�~�s�(�W8sҙ�9F	�wt�;z��m�p�|�W�h��Ϯ����滿:��;�<����G�e��Bk���O��mV���!*��]hJ���U�.���̈҂=Z�ZԁEVhB���g�e�0�Gb���V�jC��Wq��A�$�����t�CަEϷ�<��#�h@l��F����A)�P�5����)��9��̷�cí���2$S�h3�����Q� e�)=�=�D�QY� �s�!�a�~�CX��ǣ�5 �(�������vƞ!j;���%���4=e����3�^M��j�vfʓ� ���[�˟���u�r�^��B#�\�:|*�ɣ��[���)���RVޕ��o�F�W`x5�K��h4�n�8fQ���=�.�L��y�>��Y!u���3���p��UXG��d�Y�_UI�5/Si�&
Ћ�j3�z������xT��S���[�0����!�L��P>��p�ER�4�{ޣB�.��*n6ŏ6J��\��#[��g�8����G��^�ޅsrF,it����������{?�7�$���x����^;:��K���|��{>�j�Oy?���E&ݴd��RC^��u���2���46 �E�]x�9r�t�C-5�d`���'����˷c�(� *�+�pUġM�#_��^#>�mc�+n�/��"�׀�n�8�%�M��!�V�b@�878#��8���L���p���m{A�\���6���SF�UDթ���5�#U/1,��$�3�F� �B���K�$a��K�(��5������(�ȦG�wPPt<~ky�N\z�R�Ad|n�=����c#����U7� ����㡔��۶O�<E���g#`�E�B�W��	8��>�р�ãԅ	��kd�&�� ��+/�Z���ni�(4�K��o��S�����U������L���
G��Q��.���(�����Te�;��/����6�Ⴑ9֡D�[#��J�)�i�߹p]RN�f8�,�N��^j�x��x؞���������W�Eo�{�=t��������W���;�ӧ��0�#L�����&�R�Q�d}�!*Daa.�P&+��p0"Bet�$��r@8׵_��/.�xs�ݟ�a�ߊa꧈-�v�!�r~���:��L*���ar<���!�r�`*��Y���2�f��~)"�z%5���s)�XSE��s�8�,��?aВ#���;�4�j�Tzk�8Ĝ��sI�Uv�u�_�_W��3����WPM��,Ս�P�Z
ߌٛ����v�(�F2533%9s�%p�iD੏,�x@�zoJy*j&1Ӷ��5�P3(�ө��*�M�ȫ7!�&\\3ȑ��+�nRQ�B��R�5�eqH[�4��+1�c��ܜ������3���9�" ���!�m����iiC��`��Y�lA ��=�r��3R�j���H��&����*S����S�gG�����E���S�S�Ig�f�kj�YA�F��^�� v��<+^gn/��hg�l��[�x������7��+h���蛳�}�{��ƽ����/��|�= =|�b-� q�q�%�[��PR��J���T�w��~�
�/�i�����y��螐����(<�����D��#B/��� d��mN�RXnH@u�ig��mn	�׺&���G���	�����;��L.�R3d���ƭ���'<�S 3�wVO�ԛ[��L��,��r[���g�t��=�J�`�o[��w�i4��4#$�"�����������;�Tu����ic��pk���3 ����>�Lw�C9<#H~��cb��^��5�kǱ�1y�Ȅ���z,I�)����.q{�P$���օq�?K�f��8BRH'�	�9x��끘�Jը�Ayg�t�Px|��Y�g�B諢�YP�]�C�w0ė���@���]p�~��n��3��u>�h���e���O�FxM�(�w��x�q^5��W����.��[>�5��68��	�ܛb�r��C)K^@���ǃX���e���p�h'S�іx}^:I�7��� �#��>p@�3�=�n�Ҿ��/���?���I��ڷ0�\��� z����ߝ���vq�z����~�v?mG����c�ֱ6�A�qs����upp�67���?m��U�9@���oosR6A3υ���Wy�)@)���� J���F�.�b8����)=�;�	.���o��
����Q[c{�
���h/���}�^^o�K�����fi\��$����[eL��zsbkm�C{U|�x_}�p֮P�U�i3�N$�-C�S�O0�����?Fa���x�m�.�;�m��CL��z�g���2�{��j��E��BCǕ1�S�˴�A��M�{�9kgV<���ɔ='���*y�B���,�vOs�=�gw!����^[ �ǟ=��f[g��r��������(�4�<��`�	��7_��8漄���C=�Kms�~[^��)��I���Cx/���vm_����}�{����ObXV8�hoo���ڛm�Ν��`�t�v����˔���ûﾏA�l/�>��W��k�[��ýC���^6���yg��7��X�}��ez0LÍ�g��򱱱A���	�'�3��;`>y�����~����� �AP^M�ۃ_��V�֠�i����f�����������o�-Ε��1.���@c���_}%��{�-j/�>��q���mO?{�^y��6����j�����W۟��w�ڻo�����������}=����|�<����ݶ}�n{����z2�Ww�'?FI��aFv*����r�u9�+k;�y��o-�l��h�3�"r�~�@ԭ����Y��{����w�6����������)A��P����=}�E{�7 x�mol�h~T �o`Me|�œ6!���g�?owC�>9,���s���y=����!J�iW��dK��k��E��W�*��x:�����o�0i� �����־��~����ţ�|���M`닇�E)^�u�����Z'��x�I����=ϗ	M��DO:�>~�}�g�U�i���ԓ��s��}�a�|��^<l�;�����������g���y�}��'m�Uh�q8ƭ�Fu��]]�CN���c �O۽W_k�������MBk�g�s�s��+��?jo��Vh|���m~ݠ�̳�Q��(��
�n��z���AY_�G�hG���Mz�]�`�}�������T; '��ۇ�!p����6���Q8f�Xb����el`4����ѧ�+�}9��O��y)�*�TXn~������<n{tdh[����#x�����nllQ/��J���lm���{��3��{<�d�a`��E'=O�x�=y�8/=�L�r��FƽN�*g��n�����g^�D�z�E�~x�o�`��"���xEʴ/Rҋ�C����:�a�s��	���:����ڌ�vvŗ۱��3�	���oem�Ӣtd�x.;�g��&�	|"ր��(/�	�|���� 條V�$�ht
���i����}8y�;̤�����ob���{z2��	a�D�	Qy��]W_�%b_k�{��.��q������;����d��!������k��J��X#,���A�x�����㶺������	Vn���ң�#d.����:�ءIz3�;wJ�j/�yﵶ��yۄ�/��:���X	�n|mr�mfba�g�g�ݯ|�V��`p��p�����S���:�����x�7t�w<�o�c̉�o��b�����3�҂����a���JO��j'Ե���e�'M1�P����ąe5c�I�_�jr��3*3z(`��}zI<
z�v�s���s�1����70O��oFۂ��?}��,�sn��r!g�ON~��z��{�ũ��`^�
�tW5<���^�<D�`?�����vZ�g^E���%4uD�0e�һ���9 �=��d=����}��!k�^�����s�/��G��3g$NN���(Oo�!����O��LW���i�+��N�.�9�AS�7�4f�?�,�ÒE��ƈ��9"`�ٓ����W0���F�Qdד��B ��(?&���2��G�K#�\�ͽ9���3�.�Ű}��)K�&����/��4���Ϗ%P��t����a�I{�7ڌ��W�p�q�O��Ia�9
����ǁ��n��.j$t�F�(��	��*�>�m��k�����2<���C���J��:.^��*��5�L(��G	ܹe}F��T���)[Ƞ�k34�6�D�M_e���SH�(Մ�*m��(�F�}��!�r��N���==5���&��s2�gu}�a���`L�o[N]jlL�6ӛB�j%!U���ם�yn��ٙn<3&P@�O�.Ԡk�Ny|����CJ�@\��P8�@��B���űx���h�Gf:o���]'�С-�b�a�>I9�TH'D��%�@���*�M��9P����K�+h Cq�Y������1���� /mO�����;��>����&e���`�?�"�烱��������j_³��o��K]�h��d|��Ç��_�g�MZ�ᅬn�Fφ� �x�P�<ܖFw�S�%�"(���+�;J!�v�M��vw	�2�}�;k��mnm�1�b#�
�?���k[�������)��¸����DV�m)SV
ð����=��e>�H�%yI�p9h�(���������/h�N���'r���ɇ�l1�C�S:W�`lKcB8�inbN湡	�&�ڕ��0��:�݅�����]��C��V�p�q�Qm�2���~�gt����Cu�DyN5�&˜�� ����Z��Mxi��h�0�=Э_�>
����H�|��a�w1�����H�`���^0e�З�^�W�a+<��y�	�Eg��u�@g� �Cc�L�����&E$�tt�[��$r�����F�2(	��W��>�����=�{B���i �a��Ȍ����V�c��`#�W�g�߾�`����|���ĝz��0�͍��>.��L����w�p��}ǧ����K.6�L6���~۟��N�W[�=����2Mu@����v�̔.�����1���Cy1ܝ�%H,Nz�Ų��s8��*���C�_O�~N����S`��#�o���W��8߿̐Ğ��ӧ�Q�ghw��C�q��;$K�e���1(��p	��p���:�x}��5�tFp���x����^B���g#����ָ�������w�O���
A�Khx�l��l�K/`}�x{�W�Wݼ�98{r�pƉ{�1�/��OgdJl�	C�����&������8��y��/Jz����l�o~����-9�Dzd�3�{q��9f���!,/^��~��v|q�<��[݀�i ����e�6n�>�@�`��y�q{�ν-�ˏg��4Sb��O����Eb/1���50���'�v�1������Q6|�<8l��n[��@�Q f>�����U�I�Ի�������͕��O>h����O�g��������O`�ʳ�m�^e�؀cm{̛EB\"�v|}'�	AHǻG�3��8"p�s����qƹFč?��Q��`|��O��Oڹ��`_�h�P���r��ߠ���F����O�-�f+��G��P����!���ƃ� �A09cqN*M42t�1\G����H��ѫy��%q�0Ǟ�}zja<���u�=���v�!��5���*X-RC�o ����߲��2z]�)C��Ӛ3�9�K�Y�n<gH���v��Y����D�M1xK�0��r��}�����n����[`��A�g��\��V8]�-m\�`�!�I�D�-��2��(��#�p琩��%��m��mc�~\�����ߺ��?�v���5�X�Fu�:k@��K���^��x�1C�yƜ�@1P�ϣ����;-��@�eA�+7fo~���::&O�r�#�q�	��	��m��G��~�i;ssBfHq��0 �� �.�^gZ�-��kD��]]���{ī��=�;5>q�0g�~g+k`��2qÝ���21hN�b \�a�{��Κ����m�*j�v���.F�5#�8^���)��f8���c��kV1Pt�(�*�(��R1�0c�r]1�{�&�0��`;&�L]�S;�"NS��gM�
Gن�7�1�+�0����Y���F^X&̈�<�GxH.�6(;e��X�3X[ws�6`Cp�G�}x-\b��0���dAKT�N1xzU�&�=�=�	F@æ�c N�͑������������;�_����/�Dz笳ߝ\�g�,'��g���5�G;v!�r���x!ʈ�	<u����s@�(�h��vy��!^>�F.��?J���5�疷�/���lާW\�me��<A��0�&�vp�����a{�Z�1s�UN1α/��f�Ö��I7��/s<�g�`'���"��"ӂ��K|_�*�m/�O�>D�7��k[m�b��m���w��3�(�>��&S�'�!=��!�Ԙ�;h��1�8�<U�q*�3/��X\4����=%�6Ѹ��E��#shw��\���C��<�0.������3����8@���n���ޙ�u]w�4�@c� 	��HJ�HJ�,��dɉl��r�;��J�$�)���̔]S*g��x�3Sg*5I%q\r\�7yӾP�Z�I��F�h������~�uS��ΔÚK>�~���s�=�]Eױ����7��+��@�).M88K_�� ��~���[ƌ-&�K>i��"`�X��JY��vt5��k'�AQ'5��B�vD�aZ��qΦQhN ڥZ�k|�(A�C3��y�o��_��X:�z5V�.V�d�{�@���AM�]qD�p$�)q.2��P2��R��rC!q��۷Ȁ�V3#�1���27ºr�`��Ok��ʻ`R�1�O�4K�G>F.�P:�rR����4���A-JR�QI���ј�@�6��/ߚv���4�*N ߆%̪ͬ@ :��T�;ֈ.!���F�"�/@R�J8�Ʀvx�n��M��{�-� ho�c��C6���s|ù3������F�&a��q�ZfV_��I��R�u �ARa�o����䁬6JO _
q%tRK]�bp51|vU�؁�Z�����㘯[b�!<�x�����X�.����kB1;��w��L3K/b�-��D8��HVP�1� �b����3D�2|���� hJ��Ԓ�w�&�c�^��ua�?�1��(�K(�l1�`�#W���S�mѐ5Ý�� ��	��.��]�v�If�נTD�:��gܔM!.��k��e���8���[>���-���I D|Y;8��k��m+��PNO�	��:Ӑr>@D�D ���2��<%�,�\��Hp��[lw�V}�,��C�Ղ�!_��H�6oj����koQ�O� B �M�����`�U?�m
��_/�'��*��O)��"�R���|�ۻ펪6���oYSm�??1=i�Z�z���fO_8eC��6�?`խM��m�+��1Y����Z�����L)=�73����2�#O��\��c��S�l��f�Ģ}`�v��.-"�LL&!�kl��J����ѳgO��Ҵ]F�����.C��Qd�#�j%�����C@t�7�or +���ʯ1��,˔(��� p�o�>}���� ���w��ْ�{��;�Q���۷��{�͞?�4����I���WŖz�VS�L�::胆,�h4�k��mEĄ3ܤc5^{�7��Wή�rCq����8ȩ'��X4��tGBa�|�u,����3p���Z��'�}�f�( V�l��k�R�o��=�/ʄ���[���iI��% ��v�8R��������������,m��q,#� �(�b#D�D�T�
}G�x�@MP\��Ӊ)�o��F�P��=��l�[�Hڳ�{���չ���vml��_49>i�� ����W쩋W���OX�'�@3��*��!��7 ������8ǃ�ټ�Y�z>g�C3��G���
���l�=��%Q�w�	�cK�ݼs��g����ņ�:}��O�sl���C������(g˘�=�
�q�d�Bn���o�|�@�:q}��὇�;�lb�:_��YD�H)�ʙ���޽\��^�VT�,͇��C�Ѷò�3�b�iL��͛���kBѸ��P"a������rm���&6MFp��ҙ8�>�v8�/��Ag�^��mٿ�ǘ(}0��% ��#.+�qgQ\i�hrN��X�&#=�.��`�oj�]�#%��#w���۸Ϟ~���%*���[[�YQ]}fS��TII��K��c}=�J�q�ࡻ,��6[�܌��E����޼n}�گ"�>@�}�4� G��5�N�m@���}k����=����eZ7���l�f$Z�$~��t�|.����y�oVD�w.�B�v���^y{�%+�Be���*�A
>�+�C���(!G"e�L�4@��"aI����}���v�����3����1%��w55=_�!̽.9�y�HQrOq<�%�C}:O]�;t�%~�/�Mb���3�z1�O���87OR�}��2�N0�0V�e\s�Q���}��k�]��^>�q�۷�濩mh}O��d6��t���u�歍55���?15��56춣%�ƻ^�������"���"�� P
0U���HšH��n�>���6j�Q��s(AE�`	��,7$�(�0 ��#��?�4��K�ED$��!�i��������]�F"��V�d/����k�h�׎���ߘ>r�?%p���$�:������'q�l���4����n��z�^삕O[{.҈&Kp%Rn�h!�R[�+b.��&rc/E��J�okl�2t�?|�i럛|������#�?Σ�v�5�兞��mkn�8n���u2vtߝp���p����0F�I�Z��&d���H�`ՊQ�> �����'�E�*{陟���������������:y>':�7y���ؗz������am;������m��_��e&HyVCycACFi4&t�dE�~j�r�tɐ`u(��v��=v��w��Ȃ�|��DMK�}����WSSSbm����;;;_�ƣ�ܳg�__L�۪���*j�|��6��4Y��+�v�.� SK�p4����lj��d���J{��ɼ�ϻǥ��k�@�E�hwc(�&{!�`S��8��a��R�������Bp��{(�������]���힃�۹��l�}��]\�P�� �Ꟍ��}<N��鱁G��fPr��x3$�ہWj������ι𫰧 �F�!����1f�7�d��v���?����#	�u��1��3�|����M׷n�jv�2t�֔�^X��cSV��3�eF@�&E�}�B�C��]����YMᔲ��[������tҺFǳ�}೷�z���N�tk�<�^�<���Ou]����v慠�7Y#�殝ۭs��x|O�I�5�GD�qg%?�p��`P�⣂n�n)g7���w��t�O~�u)V�Ŀ���w^?.kt��!�=�d�P�'�������G����n��߷l9��Mr�X
%κ傷�/p��d��2�f�%&�Y3"(��@����j�^K���k�~�v9u���wy"�`�[�YG��^�X�d��Xٯ]�}*�=X�Ik�:0�mbp��  "�IDATpl��]��dz�C��8������\Y�()*�����HE��vn�em�i��u虝0�)�'�a_��Q�Imp�����W|Z-��Dnǖ�Z��N��<|����䭈��/�cǎ�ΏO�NP�44<e-���>��,��"��_r����ޚp]�q��G�?���'�m{}J���1��߼	q(4AH�|���_�M��^��Uh�3Qv�y��-f-6��+�MqT���8I��~(8G�̙���K��bX'v�g�B�fR�ŕ�g?��/����E��\G���~�e���W-������ި:���R��;bK� ���T��C�!���a1�3�#Ӷ��Ë�k������@0 ���=8�}����=�t^�%p�i+ �w�d(c�����m��v�L�=����,�W�wӑ��^�	/e��_ ̝捕�V�Ǒ��mE~r<��$T�N�}�u�0l�M�۶e%����������w����Ҳx���/��GW#�+B�4Z~Bqmk5�<�X��3e���5[/��(��r8�8Aq���kk7���x�C{�B��������o��\��Ņq��.���v+�[���6�w$ᕼ�b!3B��Z�j�
6��(�D$�x��g�Z�|jC����o�
������ОLb���s+sZo�Sq1:�XX�EZ#
Ȼ3Wu�`B$��KI�B�h���@",��P���
�/�Ofc���ܐB:E
��I���=�fb�Z�0x��q���¦�O�ټ  ��W�`"Ë2VB��ks�ֿe���h�N�����Bu��h�f�9ʀ�9�����ڒ�;��)kf�����%9�����/	�]�*���N�T�e�ݫ��%3��\�����b�T���LcAXX{ �
�!1�صŅ��*+�'�m#x_�������>S,i���r�ա�-A��(����D9�
Y�Ԧ%(����]a�dZ_ZXz��G}�q�n�j�9A��S���Y%1N�1dW�"�A�ᤴ�;���Ʃ�(7�,��k��<}
�6�1<y��ZJp��g�g�!	��!��#fD!�o��6�&۳ ]��G;����1{]�\�9����1f�L���6�J�W�~ѡE�7�x�r��n�o�0J�=EJ�������4+O�h5!�+ ��HVM�(�@�D�6�6������AӮA�=�ܳ82r�5�|�u:
��3��E\l�ݷ�$�k�;#�;b��0�ND+k���i�O�%&��)��-g������P?�lˊ)ь��Ke(�;E���J��i�O��_d�݊�{uD8/>rjm;�-�Y��=�77�jXY�����V��{! ����.�CЋ���m�0(�&�\W�	�\�Ћ�,{�M~�VX�z-���,7 ;*n�A7�T��*óQ;"B�0�fйf�.�T嚹�9@2�f�":�.�
�!��/X��,�b/˒KA2%�.��Z��8isV�J�@�V�LLQ2ݡ8�ٓ}�M���c݈�$^��h���Y��	`�'��������3E��@[�9<
�y����7�� �;�Xx5�a��\oO~:���4�I*䇘K�RR\!��B�V!��L�

��JS���8qB=��% ����D��*K!i`O���tC��'ۡ�g .@���J��0o���48�l83�c���Z<�[6�M���<�����l����$>D�w�>�LD���q����2`݋Oa��=����r�"wc���h{�/w(������X��"�HEp�bL��8ic�
�bQܒ�{ |J�WQE^��Զ��nZ��/~14?�.��>.A��<DZ�F
J4��?��L�MYNQ��Y z����,�OC�
���X��b�������%�y�L����W���(9��-e���ўM�,8�ʮ%�DR��E�j�I{d�xc������|i�vʽ[Y�\��u���绕D���T	8�5>��ZMHZ�S�u��^��+~I�;dRW�I�P��z-�8x��o�.�2�q���	B���h�\�s��=�~~��{�����[Ȩ�Ic�f�ѐ������[����vI^���a<2�Ƈ��$.DH��m�����1U�{�ry X��9XiI�J>��}���j񛕵�%a����
��aI�~.V���7���5��>��89���ޯЇ3x�.��]-y���A�>,��ӅSo��������N�	�k��Q@�W!N�c����Fy�*���}D{��jw���0j�q�.?�=н��������m�6)(�):�K�ܤ=�?�%A
G��P/���ةα��ʫ��T
��o��JA����wǯ��5h`�����Q@UP�7�K,�o�� H=W@�U�!��`��ʥ�`s]��?s��A~�7��玄���������E ���68=�W$IFh��H�v�ml����v3���/M����Y���P0f2<����\�os�����}��ւ�Ss� %9��O1�	U���&�W���x��π���W���g��/���%Jk���ɓ�Vч�hlm���I�� �4i+�R����{���^x���^
}��/�2�VU�+���;~�������㪹�����n�	�'�6���)b`�����H�d��(��h��vx��VQ���Ace�!yU
FU\\���NK�i�~�f���2����T�QE��'a6��uָ�O�72�zF�2H!��N&<�wSc��u_:r�ҹ�>�{<x!w�Yqx���|�b�_l��U�l�#ӣ���[����/�d��:�k(l�MQ��6�Y��P�(��n)9�J�cW��j|���?��W�e��?:|�����������@ �� ȁ�Q �o6�Y�:�f�	��Y��y��D��H�fnf�˯��������>)�,�}��w=r�h�F��l��� ���Y�qNĂqZ����'6e�v7li�0�s(}!��>��gz{{��޾/�p�s$�=��9�z�Z_��FpŚ�LkfH�SNK����R��|x��v���$.���^9\)7�+������$J�!�;i�ł�i�Y%(��ȯPq���I��oB�D��2�t���2#)J���ǐݼwљ�����Wbw�:�i5x���˗��N��z�����d�ͱ�:�)���m07c=+��
Pi�Ģ�����\,�0z#������l���!������[�y������v���������������#|����v����� �Ո/d�a6����$�-B���}�ӑi��Q�A�����I���Psl������{ro�'����K?��gN�=�؁�oňn}��;7z�f�6B�)c��1%��a��BLp�`.TҜ4��\էj�{�� B������(-)ڿo�_�;��?饧:D��J���?�>�iz|����loi���Cg���Y�z;@*RV�`| Fr�q��F3�����U4�p�fύ�I�E�[��^K��k�~�v}��;�/M2`�+b��b��g*"j��px-j� t�� ���C�� P��58pV0�o���Ī}������f�,+\��j�bj%����_�����6lN'fF+�U��p���O:_~d<�,��އ@����z���^�޺E��7W��� ����DD��e�e6��<��Wn��?�1>3���Sp$�#�=���YV���jj���l��X[�h��ܹ{�f����u�o�W�CϽ����X�|+�߷5��df4E/�#�����M��!�Y��i��X���[#�Bߵ���{�ݳe�%��p�Z w��rrf�ɡ���H�Z��x��F"��C�w����;�w[CK��bw�����"���%R�M�ta�#}�ś4>�E(x��(צ�tcܲDp���t���u�}��{m�Ԧ�H+g���MNMO}'S�{V�SYY�JB�&R��������xK]c������UX�b�a�Y,g}(�g�{�f!��?�_���({Y��/*�^ȦT�"4�p6?��{���BSQ�-�aj�ok�X���sտ���?���
�4�dA&e�ote�B,��v�	�:����-�6}6z�������{r6�?dm��b�>����Lbxdfu~$+���F3���]`ݏ�=��o��̴���s3�-����jm�v	�E�{� � ��D��|E�$��%���z/�}�pXm݉n�ֱckiQ��f�g˦VGGz�'�Vrӳ�5�H��Ё�������'	�>g�}-vAٔ诔��i�V�{q����܏����<��c�p0/gY��5�{�{�c�N;{���2�����d�S��s,ēJe'�z��K ʞ;>`!�����F�.X�F���؆H;GV�L�wAV��3D�D�)�-g�kx��I2���g���8�rs�۷�g�Ġ�1�jm�����eG��X�>]���JA���eh�.�����9�I�hu�������������¨�	;��;M,�)�N���U �<��J�S�A+|��|�zm�/ٮ�>��/���`"�*j/�R4���C�������438��<��͟��j�ī,g�@Z7%g}Ͼ�VC2�əyOb����m��]�U��v�D��6;M��N�`=��iN�ܦj��`|Q��v���� �`"+&]�֣H1��w��ږ�����X��qej�[$stC�5)� |be�5��H�Й+]v��"ђ G;�����U�4H�� dg��f�2��-[�Y[�d�W�"�a�D��葳�>V�jn%��v'��$��
ؑ(�)YC0WR�����.{��	�H�[�:K4���,�c�,z �r[�x`6��0B"P�qZb�i��V*KdI������p�<p�������E��b�c��Y!�<�f:9�c�,G����zj#v�8	���A"�L�A�S�l�Y\�Ʃb&�� �z�	��a���XX)����;qS�?�����V�/��W��V�*ģ܁�N ����&j?��h��s����P�\�`��ퟄum�����Ms�H�����Fzm���	��j!�쾝<u��{�E9jE�6Y�����8� �����zL�w�ya��Q��*K��Á���䈞�.X�ķ�H�N����;�g��s���CR[���a����$V�	Jա�h��K(�F����VH�e�U]�~Q�{�0A:�(8��B�~T������=An��&/�����D�m�c*[	:G?0K̹O?�C��K^%G�մ`���'V�m�a��|��{�Ɓ�0s3~�t�h����_C�󙗾�yR�)˖��<������dQ��v������T�����ب]�8gc��&�p��+xE6�X�~���欋E��s��4ƒzpIZ�G�HmL:�S�Ǆ}���_rؑǧ�D�(N$�"�>@W�e����rC�a���U@��u �"�P��`|x�q���ɗR�{�C�`��� ҍ���!R��Gv�j�;ɭ�ZnS�	V����������V���#���*��&%�dE��+(Zm�L���K�$ #K�L>	�EHZ{�d�W������zi� �}�u�A�`�J�l���ٌ��M0{�^�
3=�*���8F�y���GR�z�ʸk ����S����]Ă�w_����'�f���Xͦz��d[̦@���*�h%�=c�4i�EeF!H)�Drn��}I�.�YA���T#i�#���D�:��[��(�cS �����	yg7��$�9���2�QH�<y2���֏���%֦W�7�
�xy���	����W����}C@��]�q���w�N�f��R��g���JZ�^�>�+_��DIy�Τ&���RK��ۮb� ���t��"��B*��3���!8���i��R(@��-����(�Fl�[�8@��Fmfz�Ɠ	�H�hL����P�-���+����n�}D�6-rJ�n�?�p�
�|�_�G�sJ	Ҥ�#q��­(Nd5��: �L��qw�Tt�iQ�B�7�0�Ytd�� Q��#�����E�V�A%Q-!���8�����
���ԕy�('�pJx���EV�U�V�ՅUB��\!g�Y��H����t��̦�[�Vi=��"���81	G�%���#��T�����8�$C ��N�C��_��!���JX����T sD|�3QZ�"�X$s�ꫪ���L�!M��k|�8Ĵ��8����QT��iG�o�x���
;���T�I�����<"Y�Z������h�^{�XA��ܐ�֮,E5��(� �S�iUٟ3�7���kf�y�* ��1P�����rh���v��bDŝ�? �`���65?hq�O�ɍ8�,#6��&{t�M�o`E��	FZ�S/��R�-R���Y�+ �����8�p�^��VBW@�Z&g"��
���1Kk�at$�(��0cA4�cT��H$I
~S X�b�|3K.#���84s&�5��f�]�ă��ע�z�*z�$���x��ތ��5¬^�l�P�yw̖��4O�jh'|1�0"J�%
\Y,N@�����&F�B�+4�b	ZK ��W�^�5GK�6NNX)��#�͙�bИlS��k�Ģ�q�;��f+��Y���'��a��ѲyC4鱜�bp

0 �E�8�^��	���e�~�X�`��� ��ZnHQ��X�E�цH㮴`�*�Z��~���,�1�y�).����sb��&��/V�AX�Z`��F��L�.�<Z�!�^O= ��s��4��0s`[�]ȳ�"���͌ꐯ?���,�� D�8!��	i�Y��� ��$:q"G�f���U� ̔%�'D����4Wa�(�,�"94�6�1+M �4���v�0���ԑ��7w��gҼ��� U�O�����V�����$���F_�p+k5�Ħ蛽G;a���p$�S�;ɝ���t�V��֡Н25j(ì��f�]��o��C:s!�:�f|b�;���/���j��3�z���ŻC�����6{�	� �-������h�~E ���Z�=���NP���ZnH�ըR��Z?R:!��T
.|��T'���fH���d�4����A�5��5!TD�UDd �e	� �����w�!Vm����bUUO`��0���~�y{h�^�Z��H��z��,�C�!X���zX�X!��#��-ȟ�-r*S���
$�
u�E����I��S�W�8���NW���텾�t�v�z����� m�>���ԧ/�1��~?z�@�ȷ���}?�/���U�hŸ �9������ ��NT�#�ڡ�u�Q`4������Nt�"�-qK�Әx��G��+U�
��,q�09�� �n	c���@L�8#_#�."f�t;)*�<��#@	��d��� !G�`����>��% �A�g6ƂQ(.���S@�l%3�~󌈑���ᓙQ��q�k/@ ���h�qM>8p��z�����>��sN�F13cω�gtH	�����������/K���+��)�����+F�@m��"���^��@�;�=h��g(22��I"����@x��=:�>"�ʁO+_8`�u'�=�����E���ES���@u��a�����o��m�X��M�+h�ꄋ�$"�ޥ�~��CG�����uO�����I  ���G=g�(���0>k5�U�Xi���C�� �W�)������A�1�׊�1[x�N @����|�2�kE�}�fw'�d�!�#~��׳=�R��-�5�o8�/�\k��8`�=�&����,Iz`-̘�~���>ߪ��0���ߚ�ݦ��q&�\x�֚�!(���Y1�~N88��#�^_�����T�@"
?��oMq�c�fsǚ[B|�]���Yܞ����!�&�|)��r�pͿ�����y�rB"�_W#x�b[*���H�1��f~7�"/%�z-��Y�������~�*TrW�P2��i�M9��?;���]���Er��|dW߫��	3��+�+�Lo��p�Y�Y
�K������O��ы�E� yݚ�� ��kj�X�|�<�<�KH^(X��_��M .�G��8��Eo���}/�
z/§�S��Y+8��8pg�)� ~ʾ���X\sV]}��ޗ���K�w��}%n)�}�VU,���L��"�wW�����q���(Ӷ���ru�J��H<�8r·�О5A�LKx���B��� �?)B���g�9qo�X�/4T���$��O6�Nx�X��R���J;\Ӗi͖gm���I �,ny��"k� S/buXN+5��? ĈZ:M�YI.�H���3t�� �/���X�<rh$�U����*1iA!���5���&�ozD:�R�"TM� Z�N�hF��e��
[Bn�F	���"q�������UK����d���QT�J�kBh���~�Q_H��U�|��׊�B���>�b5,D�J��Տ4^z	=�վ�F���<zY��{9)�N���E�R��R���SF��R\��P�;9ٵز��4��[߬�_�?�ӱw	��;�fk 6rZ�)_�8��5E��/˟��$	nG� - ��(pf�����S3�a~S�������5U�������2��    IEND�B`�PK   א�X`�/��1  �P  /   images/c6d03bb1-8982-434f-b214-1a37938b12b0.png�zwT����ke�ā�AADz���F�P�B��5�Q�T�P"��@@�@t�^BK"Aj !-�=�o�[��w�u��ho8����9g?ϳ�w����/��� h���!h�$my��V���vI�����KA4�*����8>T
�s����C�U(44T���~A�?ܸ��Der-�!ht��{簬F��١�+��
�폌�TtXjC����ѷ������o���n�щ}��M�^x�}�uWͶ�ߔ��f�Ǵ�;n�~�Q��W��z�4���xŏ�C������W^�MZEǰ�1�{^��9���Yne[7�A� &��{.���u��}[bwI=�"�<n�l�lܨv��~�i#A77o6���ɆL�1����'MR�%j�&����!�4�UF�u���a��U�(��HNU/�"4���`G��dN������z��7T���9��\Č�ق�=eOu�Z	���Rl�ƚlGXYQ)��oVu����k"qz�g9P�4��x�T�ͳ�5!�U��i����#�-s�.�	�n�#�o�P$|Ek웅ĊKoE���K�-;᫞��H���f���0V^Ϟ
���J~��d�5ۙH�^��Qɿ=�Ƕ�%��V�._�|ǽ*?ͩl���-$n)����.mY�3���j�q�0�6��Ŭ儁��HSH$����m�ȥ�Tխ�'9��U���`�J�G���
w�(S/E�4��j��,�/��ˠl�����1��P//+n@�:�TБjgP1y�q�A�m�Zhs�03S��k~ק���SM����~���)ű��ٕi�A�rr������a��Vi�Y�v�iy-L�KTD0��B ,a<g��~oBnr���`[�R�2|�vQ�%��[��f��x�ӳ�/�D]q���;3�P����̿����b���0�jy>i�N����OX%���D��5�Բ���F���SI;s��Mv�qV��.mۘ�/"�,'��ʸ�\h�.C]�����i�ײ�ͼ�P�x�|FeS���K�f��(
� T#'9��(ٚ#uΈ^M��C6��c�?��1�4b���?/��V�*�c�h����x9�Hˈ2�l�1:f�C��ժ	t.�`���8'rVs��ޱ-x�%�X�_��ZA��>x���5i��©LU�
�{}��X|�H�뾒,���%�U�K���s(�������2}����:Z�+
����*s��,
���Yl�$��F�~۹	�2��	v^׮�s�ά���;5���&�0�+"ѥ+rm�ӑ��1�^J$i��1g��1�n���i=�)�T\?�V5�ęU����(��������öfo��dG�%��mmsk�KW�dii.����N���^�5�x�$���5�Hx7Eֵ��<�w	u2YxC=�~��%���F����	��e)�I��~�w�#"[�u;[g�C��z��ZL^4��Z�V��v�w�㬚{{ Q��/��5�p��_gp�0a��9����b�4S$C2^�x'��DbNg��e�w��I<���I����n�p���ˢ��hsl�W����!o��s�����)|�OѢ�t��؛�a��ţ��U��y�>�GzEN!q��\Z1L���|�O�`$�I�BɆ�������{&T����$x�*����V�dڄ5$�M��Dko�tD��)C����!�5ʘ�@aK|�ׇݓo��.�'�񓪮j�1��6|�x�F����G[C��&e�~�]�R��R�l2��};�b{Q��d<:J��Q�}3����mk�
���8���9��<���~��������o1ϊ6C�n�2g�!E>�GsD�?u�mN�|�1;8����jc֭�p�����Kn|�{�3f�<�SD�7�J�jPZI�Sќ%h�ED�M��+똢��[���,���� t| imj��".�_�iܔ������c��㪐J/��ƻ{m%,�̉Hw`n6+�G�:�NJD�t�U}B�0��Z}#ҍ���q޹y(��!H�'s�6�L
^�zc�#���^	�n�Q'���_�+��W�kƌ��cf����,\�����p��N�[�����I���Ss�?ݵN�I�o��I�I������j#ꪸ����&�m�?�y��)g���|�|?:�+���*�/���8�6�?���J4����SS��5���x�N$V�Q��q�!���s�dǒ1%�48����t���J��0Z�PfbvD�Q����M�"bմG�2R��#R^D��+刾E�Um������uA}�I��
�~�Շ��S�u0�u������!��d�n�Q���7����x�|��r�|�ST��kO�d��pf�G����c�'F��adyH+y;]�Q���$F"���o�ܟ�Y�����ck[\;3�*x�X�d��VDVQ��mz��4����A���0����> Ph#M�h�ī����t��[�pQ}���YY�H��EN�����n�p9�l�Q�t�sݦPM'fc�)@bc�R<�@9�?x-e)^
��-e�^�)մ�{���4� ]y1����"2o�@`7���xZ��R^y����olP��_@[I�W�K�y�)ZNx�����^�W�c�(�����Ʈ�'6�Rf����.�o��
�5!�e(:J���׳��VK�;��`�;0�[�x�aҊKG�V��\p���n[����1z	���z���i����/�Vqke0�J!!⮬�r���CJ2	��QNG�E�_J��l@#��^}���C�]�k[�2����6��]隙�x_��`��$�ʿ�\G$�����X�f��I������Lq�H7�>�D9A��-�G�ٺ�g��Zi㣊�� �3�[5�P'I>�ּ-�s��ӯ'$��0�ϓ���quwg�����j|=g��!��iy�bf|�m��/#��f����M��*	�c�-�=�v�_�R�\�@�+ŧӳ#���=���Zq���#{��	o)

��YK3`G%	�<��2	�6(݋���|tߦHs=��L|��N�>9e-�M�&3���4�C_��쭪
-+���rc(�^$?�Ɵ7w��l��$�T:��{�=G����Ҁ��ŝ�Hn�@·[
_w<��]���%�65פ'��oA��1�&�.E@P��#�ed�u,sǚi4G'�����oWL���}r�Ї;w6ut��R���������T�HGC�_�g�����ltԱZ\�>�tHH�Nir���tq���gE�t���~�������/�o�hfn��~VT gj�������Q��m�����������QGY�S5�z͏b��8�흧���QȂ�/r$����|�x�%7��cR:;��O�<�o����C��jb���y��N���B'?t�Ė]]Jq�R�Ħ�`��_�?���+����b��q������;[��ߚ���*�:g��[��(EB��f���dXF�iA_mT�w�ؙ�&~,�p����	^�8a���^��뿽ɥ�X��(�;�`l�-匬�O�X�H*|�������[��~�S�b0�{�g�ϸ����%3˧��wZ�U_�ѵ��df��pE�����K��e�]c��>��N�2e~�B	��,�Z��ב�2�����쮦�K0E�3���/�D2��������/�w���>ы���˾�j֮[:^�����9�~�{f��d��������A�����wj~Y6��-�jlg�[/,���覹�<ԛ�U.��V�t��W�(ڱ�
LyP�N�����H:�`W�?Om^5=Ë�P粤U�
�JŷJ��4¥�)޶TbK饇�⏌��h��ԔR@P���w������k�[oę��R�8;��+Vѣ��?VYG,Q[���ϟ?G�]�啜CU>\��͢5��S	����LϺ��U��uz;a?�Ϩ���L�Is :j���c�SzM����`xDطXJ��J���J�\"�
�
�ʋ�C�#k��FY~��v��k4�p���ƛU�¬v]w�IVV����Wf�/��������t�ʼ;���ã�-;���|	�OXg��r��9^^�d�Ou\�6О\S�=j�.ѻ���B�ط$n�9ԫ�ѝ*���B
������H�ۙ�vmrM�k?�L����[��k�}Q2����i%�����������A����L8&�Kg�f$�4��2n^�'�\]�z��q�ODw����vd�eK��t�ҵ����l����o����)��̋I9�sM�&'�$<�����F6z�.l�|V$s�2Z����u�k[��6�u��ٳ�S"C1h�����_t��A,n����Ξ�R��Wk��<�_����r�y#m��� �:��2^GHq�ձ�y��H*9-9E���:�ʚKM�VH�J\t��N�#Cflo;<ߐ�r��Z��~3�e���i�u�C�+����a�^&��@���c���4�'������nW7hx��I�*�ek�p1�y\ޣ�Zrڥ����SW9�fy�{���#l�	�a���ʍGV�Ը�m��T��jL�O��4f����w`���4���'"���S��B%׵	�j����{���J	O��:'6�|�|*���h	̧��o�c�I}�֥1��*a=�?�#�}7=5�1���f��v���h�0��1��t�_'�5��jd[�^g����N�H%W���D�U��=�=�S6A7�\@�S^��I����X�5�u��.'\�G=���x"��w��n9�|��-j����ʫOfٝ�3Q#�l�9DW��	J�lX�����'�N��7|L���K���)5*��S��蜜����$؛�ܹ6�A'�ezx���Z�m-��z-;�&G-`�A����� ��*�Ls�M�����U�cA7߸��R8�Jyl�B��Cc̺�W�r@���/���G��FKo	�<���? ��N�E��H��E!��V�XZ���<ҏ	\Y��x<j?�n�ˠ�	A1��BZر�y���ň�	Y��<�%	)i�w؉z��B@؉)�����W	5���@�*n��@m�@t��%>pu��Z+��ɐ�����Y�G��t�Z.s�5�I�Þ�/�{%�h���ex�Y���cd��w@�$&'[E��a�*H��fyT~.P��" 3��"e׷��PE��J�eI=�{t�r��'�Z8$.����!�^��Ō4a��&"��d��if/L��h���W���8��9��݂9���0�)(�r׏��?m�v�ݲ��E��_�f԰D.�g�;E�z]��w^
�u�W�'�=0M/D���%����э�v�y5Ń�p�	�'�WVW�Y�R�GF`?�SޖLXP$|�2��%ZWO���C��6����.KKyM����[S��t�];lj�rkm������K�RX�Yʪ�oR���,���Z}�'���RO�ϕ^�I���s�;���.�ai��A�LJ�)����%��[��T��QG��z�)ޗ2�>�c�.�.El�>��;T.��=IaHlfȒX�賌\J%�|�ر2?zi���t��홨��G�����s;��ǉ����d �w��R �DDKaYʨk!R�蚋nM��q�vOI��`�IE��דR�p�X�p���)�-����B �{!<�yƯ�;#�H�aEP�tU>�{�	�i=[n,�n{�0�5��4������Ŗ�8#T���;?<�Q����{P�3h`:l�񢽓ࣝ
��"���J��W|��K����O�!g�9I�^M��s�h/�|c-սz���;"Pc�ia��x‒Zk[W��wQ�fۧ��h=� ȣ��h<���lA7ԱjF5�a�O}�x��@u=��س���@�(W}ҧ�U����?선,��a܈�^��� �J85sc6���[�*�D�nw�1�wow".CMA�q�I��'O�Վ��i��Lt
����h %��M��`���o�N��c"��;� ��:1Y0q���gtw�6X��]ǖ��ɹ���e�g���\�{������+
����2��o��,���9���z3V����VB��sf'��p�L�����b[� �U�iX��u�X�ɓ�+���Q<���O�RY����<P,�>�X�Щou���_��Ck��.KY��ڠ�sM##�X����b�?��yJ	�{`E�/��w���X�D�X�����U��w�{�ck<%4�V
K�י^-E8酿�yȾI�5@Ғ��8�]���R5&
����A -%��bK\�����|�SL���Fe��Wn�c���� �{��+v�1ɝ�2�Sz�/�X���i?>sʲ*+V�/�$*rXK]t�O8vD���X�z&;�7��!���f��.�����k��,ż�lj�\;��x0f�X�+a�{�$��Bҁ �������@	*q��ɤ�t������l�~K�r9�4��*0ˁ� ���%i9�,<���p������[�1��S���^_\21�&���a+��)�y�;��]����(�'?7�R���]��&BL�N��e���K��x�����O8]^]k5V�����U2����N:���չ�yف9k��)H|l�;�H>���%�ef�`Z���9���3�����X7G�����9]ζ�J?�X*�}|&�N�)��7�bvqq@4ڍ���ݤP�����;�j�S ~�@QUUZ�&HV�*�][��u�D_y�@f0�B���'���T�'F?_H�ZX�Y�t�\8��R���u,o��U�p���t���U�cj6���ܖ���V5�1+��C߂i�.%��%����n���E�	�t�[,�s:��'�� e۪fJ�KV�&��Z1R��T�}�Դa^�r����7����҃r�:��X�R3i*��d��vRZ
[g6�Q���5���D����޽����u����6���|�ٲ�G�Q:Z��^�����eC�7Mͱ�a�K� �� ��	x����,\]�r��/�ݪ�9��e,v�����^���R,sY/E5�<lAa�f ��@�u&G�gG,��`O '���ݍ��x��b�~2I���?Q��M}��8e����'۽�J�h�������-!f���*���ˮ�bl�����(��=}�
װN�5��r��l�ky�HHb~8���
A:O.�|+�a��I~�����&��[{��B��u.�3��j��+f<�\և�Ù���έ�G|�yWu
h)I�sO��$Өw��C����;����ѡ�{c���;'����uc�5)��Vs53������\X�y�HZ@������:!�����5v;�L�I6Y�u+�9ft�̦\s��\��잘l�*�T��>�	-���B �����#�&G��>�������v�l̮xR��ǆ����K_Ձ�}+���W�U�������@�NYQ��k�j`E�WZK�1=i��q:RN)n����H�tiJ:P�zᣑ/P�y�G7����u�ER���I�N,E�Geh�/R�~��v�����P�S���h��	����*}��Q� ��I�̉���2u�ku�O�e��6�ͫ�/���I��O���{���Ԍf�ϥ��D�$y6y�G\A0������ӧ��"b<r���^��J������aAu���8H@NZ��+���� �4��Ҥ�ZM�2�K��-���:iR�n�4v@���˽�v��*���o~�0���%б'ݽ�/�[�&�o��������}19s0�+���@YSZ@�E�7��oR��Ջ9$��L�C��f
�'2������6�vxmM�vi�4�������%�H!\sŃ�.��f�M,|B�̶y��}���ie��>�{�.�|y��yـ���
�}�.)��w���������n��ݳq����P������$
�Zᦙ�HOOWR#�Ck��ټ�Pu�]܏3m-�j�9�,��\�]>�_����4���R��(�^,4G'�>15�1��p����\�n����?�y
w��O�a���rכ�G�7��-�?n�%k��-d����L�矒��w��t��y ��� /����3>\��4�����5<������r�o���+�w_sv/�/,,$�v��w�y�\�����/z}{�`���7C�A��w��őQ��R�B����O�U5.�*m��L��N\$M}j��i5�� �k׮�GԖi<�%b?�^�����.��'LMM�Q`ʣ_��˫��K[F�yuȃ�ѡ~����1/iSK��>}�Ժ�;<Mxu�c{;-NNk��#wi���� IÏ�*���T

¶+V�������g�AѬ��N9�F�8:������դ?��&�:l�mh����k,SX�ۧ/���iɽ��7�`��r�jK�̥d;�%v�_ĩ�Pa|�?sͅRр��PTJ��:t֏�@��嵐���$z���RU)w���|�Kr]�k��1v��,"����fP��B_�mM����R��r���ɨWI��T��Vg---�_"E>�K�*{�����i��(7%��`<�{���Ҿ����x�yf�'�O�0���?r�i�:�J��_Gg�C X��-T�ڰ�:/�q���tqk~���a�E�o�˫4�u�~�����d%uV�����z\�sx� ��Pf���SeQʴ>�x��ȣ'qu
��x��iuӣ��u��yt�/Ru;��0Am�[����蝣�(&�|�Ė�zV�'�y3"qwl[������VC��^�.�|�PVy鵵k�"_�~�S�Q���dy!lg~2���A��v]}b޸��D�L��7 Rs����@a�ֈb��Y�)���o�[�o��)C��1��kT�(_o�nn�;J�'u��v<v���Nm���Y���(iDl{U�]9�-ă%	���(48����W~a	���Qתr!��ƌ�8��'��a��/�3g����QC�ݸ�Z���Á��*��<�v�ك�bǢƧ	�͉ւ�V2���f�0^!�V�w ��~�k9��վ��n!K}d��+*��C�p@���L��Y�9b��+� ���)��i9f��rv�.ʔZ�`�3�+�E��l�Jw�^E���R�}�U�)X���:���c���؀3��8�/�`��d��{'�>��b��s�E���˴��V��XB
�͏t�6`fڭ@�M�q~Fz�<���2-V����5;),��K���Z^z��	�sj߱h�Tܝ��P�(����\���$�4x�}F�L�t8����=b*�޿Ֆw�����H��+'''u���à+3++ѥ�-�%��%w�{�'x�V���6<z�r!H={���~���#hgyo03�L-���@��������*�	5_3���:��dL h�O�Ȫ'R"�} g�*(lY5;u��L?m�`z�ժ�N����(<�<�i��XϮ��a��6���^q#�c���,u.E��A����R����;? 	y��sCS��v���k��ʾ��-�Z���9�RNHH���8t�;�G��0�2�^DzBJS��t�k�/��������GX�M�¡Y�ʡ�ȭ�=�E���:����h8���6��>�Z��l~5r(�~@���z(�/��HMi �j���K��̕3�c�w�O�TK�Ǻ�v冗���RPaNmS0��sr6���1��Ws��X����|Z�b��<8c�3B�@�^��M޿Ȥ�R/dG�Ǭ�?9�ә3M��hl�� �or��,���T;���|>�x�"\�\��C!Y�U�l-2����_|{������s'���.��`��*)ͮE�����~;w2xHp�d%!"!{�(�j����DZVا��h��ﶤ�X�-*��������U�a�t#��8�ؤ�ac��A���M��;����?b�P���k��{�2�O�c��J���P�.S�#:�Ԍ�XL���X�^`�]̈���~X�V����M�7=��3QD�Ejǌ�����������Ld�q�C0�D3�ٛ���!I�^薁��9  ��U�2�%pN1�o{~�1�K&�$d��k�m^]�����<Cty�����N������CX^܀!Z����%d�	X�e����4����@��9�S�@��I��7�y岄x�Y�p-��XC�-5ԩ�6r�����zf�3p? CF��G�&�������t�����6 ݳ�a�����/%Le�7����C��D^.�w�9�P����q-a�����+��Y9�\�+�뛱0#6$��M����f�L$� �h�0(��I��g�I� gdU9`���6�3�3�T�}�6�i�z�����YE?j��,���x�I�����N��y 0�	5�K�VaQV�ʠ�(�XRu~Nzhw|���Vlt2�b�J��o:�N�uБlI��s*Ɣ�?_<i�*bn!�2�d"����X�K�m-O>��1PPk��/? W��|�d����ڮ��Y�92)��lڿ{ҿG0��	',5�6{c��vO���\b_�KYf���DN�� ��S�fQ^����oVf<�II$� �T�bK(|��#���sY�¦P[R�Y�*���:f'�Dz�(K��ULx��Eu8ڮ�m�	�l�r���$|.FY�ʪ�n����\_�3��3/�'�V$u�B�M*{@���Y��$`,)����0N�j�
��s;���0�S�`n:Ժ�U�ܮE}�����/~�Y�i�2�d�����I}��V��n�bq�
~�=s�&M���`� �-4�r=]*�</Mb����$�h�uNZ����;9E�]C�&��e�*F�O�]��C脻�Nt�.�Db��D.�S.��Q��k�ǧ�V��,pN0~�N�@����b�I*VBsC��ЕϏ����K� ���Xz��
��dR��L��3M?+�x`�}���׾����C�J�$dΏH`��7.0�!�^Qꤐ|nU�ݲw�L��sC9��Q�;�^�uk�3���:=�/ǝ���Z��m6Έ�|X�-H�7�$��� rg���M/
B7�>�-9;Sw�0û�=�d��HR`�/
�?
�Փ�y�B��{ǆ�R�`�x����=<����fƎ��M���3 ����[4Z���HϟM�y@K\.2q3x����Q����������F��I���EL~��5l=źl����%�I�4ԕ��U`8�z�5w��d�&��S�%Xܳ�Q79}�js�5��h��U�aI�-:y-'����܃D��g�Y�����[�"j�s�|�Gm+��nH5���;D",���9JC���h����Kp���Hm���Ǟ¬��w�mB�����c� ��4[JFrl�e8��͒@�z�r�F�\XR���ӧ��K-$t]�	�P�hiJ�l��u�jz{\)�������q1ۂ�q���c�=�5!t�Е�,���f�ұ�R"�@�"i��_3��氊p��L��Ͻ\] ��t�֧^Z���mP-`����9�a���{l�����v�_�\�~[u7F�`�خ�3�b7�������� %D��;t��xy}�j
.
��Y�.�)$�D��	�s�޳=?��ޓ��M=C�7����F�-���̯)E��)��
�j����R�Y�Z!NE��?j�-�R�����6�� S��ݰ��;1+*83OIV㉹���)�v;g��ˢ� -�`h��al���X���Ě��o~��t�,Rrè����|7B�~^L7�/KV~�YՋY|^�eچ��h�[���`��������^�"���|*��V��l��R�a�W�\�mT[�A����y���ݓ=/��"Mv#�nq[�K�GӴ�Ն/u�������z���J��]ޭW�Z�_��K�6<�M��b�����>�#k�r�y����$8�f�M H%W�dns@?r��D�N�n���R���+#jX��\��� �lv �z���@}������a�X{"Iu_� 1�<0�<�7j�=�5�tr�z���|�6Qh%7,s�Z���?��/�k���c�Y�3de������-�^K<��\��s�-�M1F;P�5�t��h���p0�_�V���������}	ݜ%�R����QG4�\ON�ͷ�<�A�}�lk5ā��{`ƶT1�	�$9|�&dV��(s���	�/#��g�s����I��I|���y��p��+T;�O6.v�g�IۑC_w�8_�p��sM�$��ݻ7���4!����Mv�\;�_"8������f7��d�)��+�����NIJ�孫�e�1�h��"i���T���F��diV2#8;�)WF��x^/����d���%*%�B��}u� �y����>�1����L�1�����%#��r	r2��������}6�_���g�CohyyY��|�.��w�b��Ws�u�kM�3�Ctʆ�EҊ&��'���L�1�i�,q���&��O�	�3����r�PK   wH]Y�{&�e  �4     jsons/user_defined.json�Z�n�:���� ���%oN�i�ɥHҞ�sPE��8R�K������7͖;�%*R̓_["�ޤ���$������W?�����>��_�|�9��c<&�d�Jʦ����?6_��M��j:���y��]�O��;4������h���4I����a�@��$��������)nn�����?�h���p9_��SS�p��vYy|�����w���*u�X���#-�B����D	���6��2W�U'BC �Zd07�kM�� &�g���t����ic�����죳��Y~��bx�c��n���vf��*f0�C=�R)
��_]��Wj�����&}�g_V0��$�Z�3��N٠Xd��lO8K����c&�,�d�I�>s輙��M|ٞ�gß�ftG�1�`g�𯮢�4��:��]\�D�Y�v���_Qx�']�?����8~G�������t]��[6���G���ϗٚ�JS������.���$I-��W�(a��3Au�a�|�Z�h��B�`�83i&�
�R�+��F55�
��D5��D3����J�F�
=V��'��fڃl���Oރl�?���}���2�_g����`���wD��Y^�L�����e�;b��"�[f��óNB�0s"Ӝ�`S�:���23# �rሽ#~c����7Im�����l�ф�g�-�d|������,�����s���t�n�ԇb�h�M�F$�Yd���(¹Qî��wA8�A�W!���R��H	ON:���1nE��p��o���b�Hb�ګk"{}w�M��uQ�}�_ON�{�"������������7lv
��6���97�y�a���_���_�w��s��"ݚ.)�>[d��o�������zu�Í���*X�\��4�����$OWep���x$H���@�i	;΃��A�<�u*|J�4/'H�~�-�Ů��8�ɽuJ!Qi�v5BXQ�b�s����Hf�3IR˭f02&�3C����O��=Й'c�����G��]�����t��Z�|!����K7W��d�i�
]S����
<|Hʛ�-j��i�*�oyR��;�
�n8���찢���X���K����*���=Sp&-��������?�;���b��J��xL׏�T���֟i����+zs�bQ��|u����"�l�.�}�#1��l=R͜�&�{�O�7�r�	�a�n�~9E���&d�fu�0�>����,[����狚\�䷫zZR�����$��)�)OA7`��D��g���ø� N��%	A�h
[5�H	G�2e�NMp�k�#I�!�!$��y�B¨�|Т�}�Dش�JF��$d���"����;3�\O����6p����G�#z�|b�H�}��}��}Z�W��"���"�>�O������lP"BG��v��H���'��W��6D"p�&�������+CSlm�H9,ל��X�,O��8ؤ~������%\jȳ��>�����~9��c�����;9&�h�?��|�� fD�Ɉj���96قǰw//�g���O��� �H�Yo���^��>j��>j>�/���,/�6/vTa}an-��f��R'Lx��8�7H2E�0)&�j^w�C�p)V�Zq-�)2"����Ğȍf�/I�`�Aگ�üH�)R#3�x]��3���������1%-�������ݣ#|�r�^�l[|�����8~��ttt�Ϻ�]"6�l�i�١=���#x���^5���y�����-���a��2�m�ت#��)N�Ow�u<NӮ,5q�8G;RtJ��1$�Ў�r�Z�G�4��RBZ+�H���I�-'h��'u�ʾB�ZQ��|Y!&u�ʾR,����ܕ}�xg/��W�U�I\xh����O�I��=yW{Zg��ɓx��u�ʞ�<��X��ێ����]���I;�+'m�lG�N.���oalG¶U���v�evp�*^G�Jȶ�RD�����Գ����wo�����A7� v�L6���k5���6���6��2\�w�U��e�����p�@�h��j�&�����_.W�|_���3�R�T� A����'H+IQ`T1Ǳ�^<�����PK
   wH]Y��l��/  ��                  cirkitFile.jsonPK
   �C]Y��<u� �� /             �/  images/12ff1f2a-9049-4881-9421-35ee34297c1c.pngPK
   �F]Yo�>��q  �q  /             ># images/2cd737db-51bc-41eb-8762-f3273c40eae5.pngPK
   �C]Yu�E88� � /             U� images/41553842-fad5-42b6-aa21-339597c45c1a.pngPK
   א�Xw�'<�  �  /             �p images/48eecc1e-62ec-410c-a9f3-e9ce63fb3255.pngPK
   �C]Y�i�4�6 �6 /             �� images/67f527dc-1a08-402e-85e7-42fb10b753e8.pngPK
   �F]Y�'���U  �U  /             �� images/79f1f6d5-8698-44f6-90ff-b688d5ed2669.pngPK
   �C]YR9��b  �%  /             � images/81a2be6c-b468-4131-a428-4eb848a41f07.pngPK
   �F]Yd��  �   /             : images/83c9e9de-0e54-4db6-8a4b-a33510724988.pngPK
   �F]YN�v4	� m� /             �Z images/91e5cd07-2a88-4b0d-9128-72e2f992e16c.pngPK
   �C]YC��cx  ��  /             � images/92d0aaf4-7c05-4843-a3a7-a4d3b320fab8.pngPK
   �F]Y	��#u } /             �� images/a63a4c90-64b6-4a83-b635-c920396f8e2c.pngPK
   �F]Yԯ�|�] n� /              images/a794cf5c-4b1a-47ff-be53-d48f5d14bb41.pngPK
   �C]Yz�� 5& ( /             �^ images/aa32f2d7-3103-4396-8365-58a51d23b1a5.pngPK
   א�X`�/��1  �P  /             x� images/c6d03bb1-8982-434f-b214-1a37938b12b0.pngPK
   wH]Y�{&�e  �4               Z� jsons/user_defined.jsonPK      �  ��   